module weightMemory1(clk,address,weights);

parameter DATA_WIDTH = 32;
parameter INPUT_NODES = 100;
parameter OUTPUT_NODES = 32;

localparam TOTAL_WEIGHT_SIZE = INPUT_NODES * OUTPUT_NODES;

input clk;
input [7:0] address;
output reg [DATA_WIDTH*OUTPUT_NODES-1:0] weights;

reg [DATA_WIDTH-1:0] memory [0:TOTAL_WEIGHT_SIZE-1];

integer i;

always @ (posedge clk) begin	
	if (address > INPUT_NODES-1 || address < 0) begin
		weights = 0;
	end else begin
		for (i = 0; i < OUTPUT_NODES; i = i + 1) begin
			weights[(OUTPUT_NODES-1-i)*DATA_WIDTH+:DATA_WIDTH] = memory[(address*OUTPUT_NODES)+i];
		end
	end
end

//memory
always@(*) begin
    memory[0] = 32'hbca08236 ;
    memory[1] = 32'hbde0c38a ;
    memory[2] = 32'h3c2aebc8 ;
    memory[3] = 32'hbe1a77de ;
    memory[4] = 32'hbcd0198a ;
    memory[5] = 32'h3d80cdda ;
    memory[6] = 32'hbe28c33b ;
    memory[7] = 32'hbd7042a0 ;
    memory[8] = 32'h3d55a9b4 ;
    memory[9] = 32'hbd0805a8 ;
    memory[10] = 32'h3c1702be ;
    memory[11] = 32'h3dc98d3f ;
    memory[12] = 32'hbe039ff0 ;
    memory[13] = 32'hbe2ef8cf ;
    memory[14] = 32'hbe031d28 ;
    memory[15] = 32'h3cc02e52 ;
    memory[16] = 32'hbcc496a1 ;
    memory[17] = 32'hbdaadfbf ;
    memory[18] = 32'hbde39e44 ;
    memory[19] = 32'hbd60baa3 ;
    memory[20] = 32'hbe35ad08 ;
    memory[21] = 32'h3e0b8f42 ;
    memory[22] = 32'hbe2ec61b ;
    memory[23] = 32'h3da802ba ;
    memory[24] = 32'hbdf8f2fa ;
    memory[25] = 32'h3d79a773 ;
    memory[26] = 32'hbe02bbb9 ;
    memory[27] = 32'hbddcc137 ;
    memory[28] = 32'h3c8fa1af ;
    memory[29] = 32'h3d6c70c9 ;
    memory[30] = 32'hbe119599 ;
    memory[31] = 32'h3cb1d563 ;
    memory[32] = 32'hbe37e736 ;
    memory[33] = 32'h3c3ce899 ;
    memory[34] = 32'hbdb5818a ;
    memory[35] = 32'h3d166dba ;
    memory[36] = 32'hbde9a069 ;
    memory[37] = 32'h3c3febe6 ;
    memory[38] = 32'h3e0a20cf ;
    memory[39] = 32'h3ce4be9b ;
    memory[40] = 32'hbe347797 ;
    memory[41] = 32'hbc2152ca ;
    memory[42] = 32'hbe0db1bd ;
    memory[43] = 32'h3d452b7e ;
    memory[44] = 32'h3c751939 ;
    memory[45] = 32'h3dc3c205 ;
    memory[46] = 32'hbdc46430 ;
    memory[47] = 32'h3e023359 ;
    memory[48] = 32'hbd8c1c8a ;
    memory[49] = 32'hbbcad94b ;
    memory[50] = 32'h3db94cf7 ;
    memory[51] = 32'h3e4529c2 ;
    memory[52] = 32'hbdc77dd1 ;
    memory[53] = 32'hbb7b81a0 ;
    memory[54] = 32'h3e0df28e ;
    memory[55] = 32'hbde6d568 ;
    memory[56] = 32'hbe130a19 ;
    memory[57] = 32'h3dfa1adc ;
    memory[58] = 32'h3d0be50f ;
    memory[59] = 32'h3dfeaa54 ;
    memory[60] = 32'hbe039c4b ;
    memory[61] = 32'hbe0a48b3 ;
    memory[62] = 32'h3e12d2e5 ;
    memory[63] = 32'h3da0610a ;
    memory[64] = 32'h3de94611 ;
    memory[65] = 32'hbde04607 ;
    memory[66] = 32'h3e0e4791 ;
    memory[67] = 32'h3e2f34de ;
    memory[68] = 32'hbdc66ccb ;
    memory[69] = 32'h3c010e6e ;
    memory[70] = 32'h3cf7ca91 ;
    memory[71] = 32'hbca60f7e ;
    memory[72] = 32'h3e11fb95 ;
    memory[73] = 32'h3dd1bfce ;
    memory[74] = 32'hbe3dfd5f ;
    memory[75] = 32'hbbcd43c7 ;
    memory[76] = 32'h3d25c832 ;
    memory[77] = 32'h3c7ca91e ;
    memory[78] = 32'h3ae10129 ;
    memory[79] = 32'hbe09d94e ;
    memory[80] = 32'hbe3aff82 ;
    memory[81] = 32'hbd66047f ;
    memory[82] = 32'h3e23a52f ;
    memory[83] = 32'hbdefe57f ;
    memory[84] = 32'h3e05cc0a ;
    memory[85] = 32'hbe22ea1f ;
    memory[86] = 32'hbd5f7b87 ;
    memory[87] = 32'hbc90be29 ;
    memory[88] = 32'hbe0d5791 ;
    memory[89] = 32'hbe4e7da5 ;
    memory[90] = 32'h3da70502 ;
    memory[91] = 32'h3da69bbf ;
    memory[92] = 32'hbe36c0a0 ;
    memory[93] = 32'h3db2258a ;
    memory[94] = 32'h3df55f2c ;
    memory[95] = 32'h3df2ac1b ;
    memory[96] = 32'h3e3e0249 ;
    memory[97] = 32'hbc1d1d14 ;
    memory[98] = 32'hbe09ad6e ;
    memory[99] = 32'hbd020c3a ;
    memory[100] = 32'h3e246d18 ;
    memory[101] = 32'h3e3494f0 ;
    memory[102] = 32'h3e1eefe7 ;
    memory[103] = 32'h3c5c2798 ;
    memory[104] = 32'hbd694718 ;
    memory[105] = 32'h3cfaa702 ;
    memory[106] = 32'hbd5aba7e ;
    memory[107] = 32'h3cfcdbce ;
    memory[108] = 32'h3c39ae4e ;
    memory[109] = 32'hbe18a1f9 ;
    memory[110] = 32'h3dc12b03 ;
    memory[111] = 32'h3c74af3f ;
    memory[112] = 32'h3cd295af ;
    memory[113] = 32'h3e2bc751 ;
    memory[114] = 32'h3c556b92 ;
    memory[115] = 32'h3df40af8 ;
    memory[116] = 32'hbe136595 ;
    memory[117] = 32'h3da773bb ;
    memory[118] = 32'hbd839a33 ;
    memory[119] = 32'h3e41f082 ;
    memory[120] = 32'hbcdb1bfa ;
    memory[121] = 32'hbe270959 ;
    memory[122] = 32'hbe2116a5 ;
    memory[123] = 32'h3d316e50 ;
    memory[124] = 32'hbe330855 ;
    memory[125] = 32'hbe11437e ;
    memory[126] = 32'h3e25c0eb ;
    memory[127] = 32'h3e36e996 ;
    memory[128] = 32'h3d932474 ;
    memory[129] = 32'h3de28bb6 ;
    memory[130] = 32'hbe266430 ;
    memory[131] = 32'h3e0ff7fa ;
    memory[132] = 32'h3ce3de2b ;
    memory[133] = 32'h3e45e1c7 ;
    memory[134] = 32'h3e0ed87b ;
    memory[135] = 32'hbd8d20ab ;
    memory[136] = 32'h3e1dc518 ;
    memory[137] = 32'hbdd60695 ;
    memory[138] = 32'hbe1abfa3 ;
    memory[139] = 32'hbdd8819b ;
    memory[140] = 32'h3dd06c45 ;
    memory[141] = 32'hbda5ae43 ;
    memory[142] = 32'hbd604d4a ;
    memory[143] = 32'hbcbd6620 ;
    memory[144] = 32'hbe0342b2 ;
    memory[145] = 32'hbd9a38ed ;
    memory[146] = 32'h3d7d0a92 ;
    memory[147] = 32'h3ddcfc73 ;
    memory[148] = 32'hbd3bc696 ;
    memory[149] = 32'hbc782d93 ;
    memory[150] = 32'hbdb350f7 ;
    memory[151] = 32'hbe215454 ;
    memory[152] = 32'hbdf59a29 ;
    memory[153] = 32'h3e1dffc7 ;
    memory[154] = 32'h3dd878cb ;
    memory[155] = 32'h3d80abb9 ;
    memory[156] = 32'h3d8342c4 ;
    memory[157] = 32'hbd8c69ac ;
    memory[158] = 32'hbd8d6314 ;
    memory[159] = 32'hbe0c8802 ;
    memory[160] = 32'hbe118f26 ;
    memory[161] = 32'hbd8606fc ;
    memory[162] = 32'hbd4882a3 ;
    memory[163] = 32'hbdcfc971 ;
    memory[164] = 32'h3d869497 ;
    memory[165] = 32'hbe15ff65 ;
    memory[166] = 32'hbde73db4 ;
    memory[167] = 32'hbe5a3da5 ;
    memory[168] = 32'hbdb0ec6f ;
    memory[169] = 32'h3c3169c4 ;
    memory[170] = 32'hbe18da42 ;
    memory[171] = 32'hbdb5f3b1 ;
    memory[172] = 32'hbe1f0d86 ;
    memory[173] = 32'h3de40297 ;
    memory[174] = 32'hbd0e1d7b ;
    memory[175] = 32'h3d05a38a ;
    memory[176] = 32'hbe1b09c4 ;
    memory[177] = 32'hbdce8e9f ;
    memory[178] = 32'h3dbc87ef ;
    memory[179] = 32'h3e3bb3b1 ;
    memory[180] = 32'hbcd91135 ;
    memory[181] = 32'h3d257895 ;
    memory[182] = 32'hbdd91399 ;
    memory[183] = 32'hbe0ac54c ;
    memory[184] = 32'hbc21fd5c ;
    memory[185] = 32'hbd7ea749 ;
    memory[186] = 32'hbd874441 ;
    memory[187] = 32'h3e1b707f ;
    memory[188] = 32'h3e12bc5c ;
    memory[189] = 32'h3dedfdbf ;
    memory[190] = 32'hbd86aaa9 ;
    memory[191] = 32'h3cc2b1fa ;
    memory[192] = 32'hbdfd2245 ;
    memory[193] = 32'h3de8fa6b ;
    memory[194] = 32'h3d4c65fc ;
    memory[195] = 32'h3d1a563c ;
    memory[196] = 32'h3d07e61c ;
    memory[197] = 32'h3da962d9 ;
    memory[198] = 32'hbdde6047 ;
    memory[199] = 32'hbd9fc3f3 ;
    memory[200] = 32'h3df6cebc ;
    memory[201] = 32'h3d5f6b47 ;
    memory[202] = 32'hbdfe7892 ;
    memory[203] = 32'hbd4c4483 ;
    memory[204] = 32'h3cdefbee ;
    memory[205] = 32'h3dfb5479 ;
    memory[206] = 32'h3e2b66fb ;
    memory[207] = 32'hbd1868ee ;
    memory[208] = 32'hbe15a51b ;
    memory[209] = 32'h3d4a279e ;
    memory[210] = 32'hbe2f8154 ;
    memory[211] = 32'hbbea19da ;
    memory[212] = 32'hbd935cd1 ;
    memory[213] = 32'h3d9f7712 ;
    memory[214] = 32'hbc6feddb ;
    memory[215] = 32'h3e22aa62 ;
    memory[216] = 32'hbe14848c ;
    memory[217] = 32'hbc79a499 ;
    memory[218] = 32'hbdd8e764 ;
    memory[219] = 32'hbcc45602 ;
    memory[220] = 32'hbb55c72e ;
    memory[221] = 32'h3d69fdd7 ;
    memory[222] = 32'h3d678d88 ;
    memory[223] = 32'hbdac3476 ;
    memory[224] = 32'hbe025a5e ;
    memory[225] = 32'h3c4d1393 ;
    memory[226] = 32'hbe2d298e ;
    memory[227] = 32'h3dfe84ce ;
    memory[228] = 32'h3deab054 ;
    memory[229] = 32'hbe0617e0 ;
    memory[230] = 32'hbde4ae6b ;
    memory[231] = 32'hbdd71934 ;
    memory[232] = 32'hbc12a24b ;
    memory[233] = 32'h3dffaeb2 ;
    memory[234] = 32'hbcb54153 ;
    memory[235] = 32'h3d04a26a ;
    memory[236] = 32'hbd85ec9a ;
    memory[237] = 32'hbdda8f7d ;
    memory[238] = 32'hbddd68c2 ;
    memory[239] = 32'hbdd390fd ;
    memory[240] = 32'h3cd69007 ;
    memory[241] = 32'hbe331e25 ;
    memory[242] = 32'hbe3095f2 ;
    memory[243] = 32'hbb9b50ff ;
    memory[244] = 32'hbd21360e ;
    memory[245] = 32'hbd4b46b0 ;
    memory[246] = 32'hbd20611b ;
    memory[247] = 32'h3d3b87ba ;
    memory[248] = 32'h3d345eda ;
    memory[249] = 32'hbdc0f657 ;
    memory[250] = 32'hbe027c90 ;
    memory[251] = 32'hbd3323a3 ;
    memory[252] = 32'hbd42abb8 ;
    memory[253] = 32'hbe4e54dc ;
    memory[254] = 32'h3e17e4b1 ;
    memory[255] = 32'h3deb55c7 ;
    memory[256] = 32'hbe22f92b ;
    memory[257] = 32'h3e4b94f7 ;
    memory[258] = 32'hbb9ef6b4 ;
    memory[259] = 32'hbc33d3c6 ;
    memory[260] = 32'h3e1b9c27 ;
    memory[261] = 32'h3e2385b8 ;
    memory[262] = 32'hbd8a4af2 ;
    memory[263] = 32'h3e595f72 ;
    memory[264] = 32'hbde2dbc8 ;
    memory[265] = 32'hbda5b147 ;
    memory[266] = 32'h3d7f6690 ;
    memory[267] = 32'hbdf177fd ;
    memory[268] = 32'h3d9b3169 ;
    memory[269] = 32'hbd8c58b7 ;
    memory[270] = 32'hbcbf2beb ;
    memory[271] = 32'hbdaaaeb4 ;
    memory[272] = 32'h3e16dc18 ;
    memory[273] = 32'hbc332e5d ;
    memory[274] = 32'h3d193565 ;
    memory[275] = 32'hbcbeddef ;
    memory[276] = 32'h3e11c11d ;
    memory[277] = 32'h3dc8c79f ;
    memory[278] = 32'hbcd04243 ;
    memory[279] = 32'h3e125d6a ;
    memory[280] = 32'h3da74117 ;
    memory[281] = 32'h3d4c32e8 ;
    memory[282] = 32'hbce50c21 ;
    memory[283] = 32'h3c3c0f2d ;
    memory[284] = 32'hbdff527b ;
    memory[285] = 32'h3ddc573f ;
    memory[286] = 32'h3e0b0dca ;
    memory[287] = 32'hbe4dc0de ;
    memory[288] = 32'h3d9de346 ;
    memory[289] = 32'hbe2b4d3a ;
    memory[290] = 32'h3cdd6693 ;
    memory[291] = 32'h3dca9f6b ;
    memory[292] = 32'h3da4147f ;
    memory[293] = 32'h3d8e38fe ;
    memory[294] = 32'h3e02a274 ;
    memory[295] = 32'hbe196c62 ;
    memory[296] = 32'hbbb8d346 ;
    memory[297] = 32'hbe12e534 ;
    memory[298] = 32'h3e2541cf ;
    memory[299] = 32'hbdd0ac96 ;
    memory[300] = 32'hbd664524 ;
    memory[301] = 32'h3d913572 ;
    memory[302] = 32'hbceb4129 ;
    memory[303] = 32'hbcbdd571 ;
    memory[304] = 32'h3e018a87 ;
    memory[305] = 32'h3dec1b88 ;
    memory[306] = 32'h3bd2da1e ;
    memory[307] = 32'h3de62400 ;
    memory[308] = 32'hbcf40062 ;
    memory[309] = 32'hbdf196a5 ;
    memory[310] = 32'h3d94a986 ;
    memory[311] = 32'h3de14f1a ;
    memory[312] = 32'hbdac2089 ;
    memory[313] = 32'h3b1f9611 ;
    memory[314] = 32'hbe19e70d ;
    memory[315] = 32'h3d7c74cb ;
    memory[316] = 32'h3dc76a68 ;
    memory[317] = 32'h3dab8de4 ;
    memory[318] = 32'hbd97f024 ;
    memory[319] = 32'hbc70e9a9 ;
    memory[320] = 32'h3cf83dc1 ;
    memory[321] = 32'hbd14816e ;
    memory[322] = 32'hbe3c79de ;
    memory[323] = 32'hbe1c28ab ;
    memory[324] = 32'hbd8c9654 ;
    memory[325] = 32'h3d2feac0 ;
    memory[326] = 32'h3cfd15de ;
    memory[327] = 32'h3e5ed3cf ;
    memory[328] = 32'hbe09c19b ;
    memory[329] = 32'hbd2c315b ;
    memory[330] = 32'h3df14ed2 ;
    memory[331] = 32'h3d9bf5f7 ;
    memory[332] = 32'hbd3eec3b ;
    memory[333] = 32'h3db496c7 ;
    memory[334] = 32'h3e292c56 ;
    memory[335] = 32'h3e24bfa7 ;
    memory[336] = 32'hbdc0b250 ;
    memory[337] = 32'h3cff8fb4 ;
    memory[338] = 32'hbe5aa3c9 ;
    memory[339] = 32'hbc7d7cab ;
    memory[340] = 32'h3e32e6da ;
    memory[341] = 32'h3d914f83 ;
    memory[342] = 32'hbdb0fc19 ;
    memory[343] = 32'h3d48e967 ;
    memory[344] = 32'h3d6c3e09 ;
    memory[345] = 32'hbc7f580a ;
    memory[346] = 32'h3e487f14 ;
    memory[347] = 32'hbe29ba27 ;
    memory[348] = 32'hbd276c38 ;
    memory[349] = 32'h3dfa9870 ;
    memory[350] = 32'h3e3adacd ;
    memory[351] = 32'h3d51fc6f ;
    memory[352] = 32'h3dce3cab ;
    memory[353] = 32'h3db8e6a6 ;
    memory[354] = 32'h3dcadc52 ;
    memory[355] = 32'hbe145dbc ;
    memory[356] = 32'hbe10cd3c ;
    memory[357] = 32'h3c9a64cb ;
    memory[358] = 32'h3e138f7b ;
    memory[359] = 32'h3e10cf19 ;
    memory[360] = 32'hbdfc29ca ;
    memory[361] = 32'hbd919ada ;
    memory[362] = 32'h3b9aac33 ;
    memory[363] = 32'hbd1089e1 ;
    memory[364] = 32'h3e24033d ;
    memory[365] = 32'h3bd4b472 ;
    memory[366] = 32'h3db56be5 ;
    memory[367] = 32'hbdd74d69 ;
    memory[368] = 32'hbdaa4d21 ;
    memory[369] = 32'h3db6508e ;
    memory[370] = 32'h3e5d1226 ;
    memory[371] = 32'h3ce420b6 ;
    memory[372] = 32'hbe07ca4e ;
    memory[373] = 32'h3c95063a ;
    memory[374] = 32'hbe447997 ;
    memory[375] = 32'hbcfebd0e ;
    memory[376] = 32'h3d66ec80 ;
    memory[377] = 32'h3db2589a ;
    memory[378] = 32'h3d03833e ;
    memory[379] = 32'h3c9c8b48 ;
    memory[380] = 32'h3d546ee7 ;
    memory[381] = 32'hbd555507 ;
    memory[382] = 32'h3e07b144 ;
    memory[383] = 32'h3e2591a5 ;
    memory[384] = 32'h3dd00faf ;
    memory[385] = 32'hbe2a1e44 ;
    memory[386] = 32'h3e33c1f8 ;
    memory[387] = 32'hbd64f14f ;
    memory[388] = 32'h3c8cbacd ;
    memory[389] = 32'h3e2c9806 ;
    memory[390] = 32'hbda183da ;
    memory[391] = 32'h3e01caff ;
    memory[392] = 32'hbe41b32b ;
    memory[393] = 32'hbe1dc10e ;
    memory[394] = 32'h3e4f5f8b ;
    memory[395] = 32'h38ad39c5 ;
    memory[396] = 32'hbe3bcc0f ;
    memory[397] = 32'hbe207fb1 ;
    memory[398] = 32'h3d103232 ;
    memory[399] = 32'hbdbb406e ;
    memory[400] = 32'h3e0ae24e ;
    memory[401] = 32'h3e0caf22 ;
    memory[402] = 32'hb9d059cd ;
    memory[403] = 32'h3e2e2f65 ;
    memory[404] = 32'h3d3db33f ;
    memory[405] = 32'h3c050230 ;
    memory[406] = 32'hbd4610f1 ;
    memory[407] = 32'hbdaba34e ;
    memory[408] = 32'h3df1d6cc ;
    memory[409] = 32'h3e24f734 ;
    memory[410] = 32'h3d736828 ;
    memory[411] = 32'h3d0b5175 ;
    memory[412] = 32'h3da5d6fe ;
    memory[413] = 32'h3e10616f ;
    memory[414] = 32'hbd5c4ddc ;
    memory[415] = 32'hbdb46a73 ;
    memory[416] = 32'hbccdc084 ;
    memory[417] = 32'h3cf6349d ;
    memory[418] = 32'h3e4d9ba7 ;
    memory[419] = 32'hbd9d90ed ;
    memory[420] = 32'h3cd2ac59 ;
    memory[421] = 32'hbe5731d0 ;
    memory[422] = 32'hbe496dc4 ;
    memory[423] = 32'hbce312be ;
    memory[424] = 32'hbdde5ae7 ;
    memory[425] = 32'h3dfc7f9e ;
    memory[426] = 32'hbd23a07b ;
    memory[427] = 32'h3e08952f ;
    memory[428] = 32'hbda71e3f ;
    memory[429] = 32'h3dc07bac ;
    memory[430] = 32'hbd277c2d ;
    memory[431] = 32'h3dd561ed ;
    memory[432] = 32'hbc1ca662 ;
    memory[433] = 32'hbe0e7330 ;
    memory[434] = 32'h3bc012af ;
    memory[435] = 32'h3dd6b9bf ;
    memory[436] = 32'h3ce84d35 ;
    memory[437] = 32'hbca9493c ;
    memory[438] = 32'h3e2ac07f ;
    memory[439] = 32'h3d54bbc3 ;
    memory[440] = 32'hbd55a1b7 ;
    memory[441] = 32'hbd43de00 ;
    memory[442] = 32'hbdfd44a9 ;
    memory[443] = 32'hbe0e1bf9 ;
    memory[444] = 32'hbe6e5bd1 ;
    memory[445] = 32'h3d5cda3c ;
    memory[446] = 32'h3d6de7bb ;
    memory[447] = 32'hbd537eb0 ;
    memory[448] = 32'h3d960339 ;
    memory[449] = 32'hbe12f89b ;
    memory[450] = 32'hbdb55fca ;
    memory[451] = 32'hbd84f135 ;
    memory[452] = 32'hbe375bef ;
    memory[453] = 32'h3dac6295 ;
    memory[454] = 32'hbd9e3239 ;
    memory[455] = 32'h3e3b9c2f ;
    memory[456] = 32'hbe290c00 ;
    memory[457] = 32'h3e3eb466 ;
    memory[458] = 32'hbd3419d6 ;
    memory[459] = 32'hbc257203 ;
    memory[460] = 32'hbe0cd800 ;
    memory[461] = 32'h3d8606de ;
    memory[462] = 32'hbc8de3d7 ;
    memory[463] = 32'h3cb40d04 ;
    memory[464] = 32'hbd053303 ;
    memory[465] = 32'h3e2e0495 ;
    memory[466] = 32'hbded5d06 ;
    memory[467] = 32'h3db6261a ;
    memory[468] = 32'h3c3b6f2a ;
    memory[469] = 32'hbc889315 ;
    memory[470] = 32'h3ba7ff32 ;
    memory[471] = 32'h3e2d9817 ;
    memory[472] = 32'hbd80a54a ;
    memory[473] = 32'hbd91b6e5 ;
    memory[474] = 32'hbda14a4a ;
    memory[475] = 32'hbcd19caa ;
    memory[476] = 32'hbe30c24e ;
    memory[477] = 32'hbcd4c80b ;
    memory[478] = 32'h3e3d97d1 ;
    memory[479] = 32'h3cdf4884 ;
    memory[480] = 32'h3db3be88 ;
    memory[481] = 32'hbd8b099c ;
    memory[482] = 32'hbd994093 ;
    memory[483] = 32'h3dd61dc8 ;
    memory[484] = 32'h3e292c53 ;
    memory[485] = 32'h3e32a15a ;
    memory[486] = 32'hbe317ac6 ;
    memory[487] = 32'hbdf04f65 ;
    memory[488] = 32'hbe1095c1 ;
    memory[489] = 32'h3e35beeb ;
    memory[490] = 32'h3d7a6ddc ;
    memory[491] = 32'h3b1aadfe ;
    memory[492] = 32'h3d9737ba ;
    memory[493] = 32'hbd945642 ;
    memory[494] = 32'hbe4a9280 ;
    memory[495] = 32'h3d9c7441 ;
    memory[496] = 32'h3e3a5624 ;
    memory[497] = 32'h3e0e15f5 ;
    memory[498] = 32'h3de9530c ;
    memory[499] = 32'h3e152742 ;
    memory[500] = 32'h3c0e6c15 ;
    memory[501] = 32'hbe15c6ea ;
    memory[502] = 32'h3bba968f ;
    memory[503] = 32'hbe453b8c ;
    memory[504] = 32'hbe282d3f ;
    memory[505] = 32'hbdced737 ;
    memory[506] = 32'hbd5b9629 ;
    memory[507] = 32'h3e0d3391 ;
    memory[508] = 32'hbdbfe97d ;
    memory[509] = 32'hbd651816 ;
    memory[510] = 32'h3e062ab8 ;
    memory[511] = 32'hbe17974b ;
    memory[512] = 32'hbb8048e8 ;
    memory[513] = 32'h3d6ecdd8 ;
    memory[514] = 32'h3e0da2cb ;
    memory[515] = 32'hbd582fe5 ;
    memory[516] = 32'hbdcd2c90 ;
    memory[517] = 32'h3d57c5b2 ;
    memory[518] = 32'h3e374fcb ;
    memory[519] = 32'hbde030f8 ;
    memory[520] = 32'hbbbf2b63 ;
    memory[521] = 32'hbcdee10e ;
    memory[522] = 32'hbe0d2fdb ;
    memory[523] = 32'h3e2276e5 ;
    memory[524] = 32'h3e0afd0b ;
    memory[525] = 32'h3decf491 ;
    memory[526] = 32'h3e0cad32 ;
    memory[527] = 32'hbd83bab2 ;
    memory[528] = 32'h3d710d4a ;
    memory[529] = 32'hbc12a7d1 ;
    memory[530] = 32'h3e0a54c3 ;
    memory[531] = 32'h3e105dd3 ;
    memory[532] = 32'h3d00aaf4 ;
    memory[533] = 32'h3d9e1b0c ;
    memory[534] = 32'h3e226c88 ;
    memory[535] = 32'h3e0dd99f ;
    memory[536] = 32'h3dce277c ;
    memory[537] = 32'hbd0903c9 ;
    memory[538] = 32'hbd95cfa2 ;
    memory[539] = 32'h3d95c7d1 ;
    memory[540] = 32'hbddb2001 ;
    memory[541] = 32'h3cb046de ;
    memory[542] = 32'hbda0fb4b ;
    memory[543] = 32'h3df98bee ;
    memory[544] = 32'h3d27af01 ;
    memory[545] = 32'h3e2582ea ;
    memory[546] = 32'h3e4862bf ;
    memory[547] = 32'hbd80d581 ;
    memory[548] = 32'h3d39bf60 ;
    memory[549] = 32'h3dfa0060 ;
    memory[550] = 32'hbd81daf5 ;
    memory[551] = 32'h3d17ac46 ;
    memory[552] = 32'h3e12248f ;
    memory[553] = 32'hbdd39b2b ;
    memory[554] = 32'hbcc2209e ;
    memory[555] = 32'h3e061320 ;
    memory[556] = 32'h3cd8c458 ;
    memory[557] = 32'h3e112b72 ;
    memory[558] = 32'hbe2b8257 ;
    memory[559] = 32'h3e4ca1e6 ;
    memory[560] = 32'hbddc7368 ;
    memory[561] = 32'hbe10625f ;
    memory[562] = 32'hbdb90ba2 ;
    memory[563] = 32'h3d56776f ;
    memory[564] = 32'hbdf2a79b ;
    memory[565] = 32'hbdd973e1 ;
    memory[566] = 32'hbd8c9918 ;
    memory[567] = 32'h3d4b6e3f ;
    memory[568] = 32'h3e1699a7 ;
    memory[569] = 32'h3e0129be ;
    memory[570] = 32'h3e1d83df ;
    memory[571] = 32'hbe0eaf7a ;
    memory[572] = 32'hbe145d07 ;
    memory[573] = 32'hbe2c7342 ;
    memory[574] = 32'hbe0940a1 ;
    memory[575] = 32'h3e1048af ;
    memory[576] = 32'h3d1305ab ;
    memory[577] = 32'hbe033f0a ;
    memory[578] = 32'h3e40f420 ;
    memory[579] = 32'h3d970cec ;
    memory[580] = 32'hbd018175 ;
    memory[581] = 32'hbd11010b ;
    memory[582] = 32'h3e02d430 ;
    memory[583] = 32'h3c72b7d4 ;
    memory[584] = 32'h3e34086e ;
    memory[585] = 32'h3d0c0c84 ;
    memory[586] = 32'hbc862b1b ;
    memory[587] = 32'h3d795792 ;
    memory[588] = 32'hbdac11fe ;
    memory[589] = 32'hbdc2a0b5 ;
    memory[590] = 32'h3c5dfdd5 ;
    memory[591] = 32'hbd939012 ;
    memory[592] = 32'h3d8b2a67 ;
    memory[593] = 32'hbdb9edc8 ;
    memory[594] = 32'h3d98c923 ;
    memory[595] = 32'h3de6a021 ;
    memory[596] = 32'hba38a712 ;
    memory[597] = 32'h3d269507 ;
    memory[598] = 32'hbd8a4095 ;
    memory[599] = 32'hbe436e0f ;
    memory[600] = 32'hbdf6596c ;
    memory[601] = 32'hbd0d290b ;
    memory[602] = 32'hbe13a605 ;
    memory[603] = 32'h3d7d6966 ;
    memory[604] = 32'hbc18a761 ;
    memory[605] = 32'h3c80e772 ;
    memory[606] = 32'h3d69529c ;
    memory[607] = 32'hbe3c14bd ;
    memory[608] = 32'h3d018c54 ;
    memory[609] = 32'hbdf0100a ;
    memory[610] = 32'h3d17e2a7 ;
    memory[611] = 32'hbe2319dc ;
    memory[612] = 32'hbe19b35a ;
    memory[613] = 32'hbdfd7850 ;
    memory[614] = 32'hbc9f64a0 ;
    memory[615] = 32'h3c8b888d ;
    memory[616] = 32'h3e4c9c08 ;
    memory[617] = 32'h3d961a42 ;
    memory[618] = 32'h3e022fa4 ;
    memory[619] = 32'hbc830431 ;
    memory[620] = 32'h3e39e851 ;
    memory[621] = 32'h3c956bcc ;
    memory[622] = 32'h3d7567ba ;
    memory[623] = 32'hbd810336 ;
    memory[624] = 32'hbe167943 ;
    memory[625] = 32'h3e068a32 ;
    memory[626] = 32'hbdbe582f ;
    memory[627] = 32'hb882fc4c ;
    memory[628] = 32'h3daf59cf ;
    memory[629] = 32'hbdfa1a7e ;
    memory[630] = 32'h3da2a2bc ;
    memory[631] = 32'hbdddf0f3 ;
    memory[632] = 32'hbdb75f7e ;
    memory[633] = 32'h3d2f047e ;
    memory[634] = 32'h3dc601ab ;
    memory[635] = 32'hbdc16b9a ;
    memory[636] = 32'h3e4abd1c ;
    memory[637] = 32'hbde42064 ;
    memory[638] = 32'h3de51780 ;
    memory[639] = 32'h3dd8a2fb ;
    memory[640] = 32'h3b58476f ;
    memory[641] = 32'h3db40885 ;
    memory[642] = 32'hbe070fad ;
    memory[643] = 32'hbdc92c57 ;
    memory[644] = 32'hbd35abde ;
    memory[645] = 32'h3e071620 ;
    memory[646] = 32'h3de8ba09 ;
    memory[647] = 32'h3dc625bd ;
    memory[648] = 32'h3d85d358 ;
    memory[649] = 32'hbd3a024c ;
    memory[650] = 32'hbe123dc3 ;
    memory[651] = 32'hbc775f6e ;
    memory[652] = 32'h3da6e843 ;
    memory[653] = 32'h3d441cfa ;
    memory[654] = 32'hbd50f8f2 ;
    memory[655] = 32'h3b9d545a ;
    memory[656] = 32'hbdea4ca2 ;
    memory[657] = 32'hbd77b2a2 ;
    memory[658] = 32'h3e03f4eb ;
    memory[659] = 32'hbe3e331e ;
    memory[660] = 32'hbe24665c ;
    memory[661] = 32'hbd7feba9 ;
    memory[662] = 32'h3e1dce8f ;
    memory[663] = 32'hbde93c09 ;
    memory[664] = 32'hbd6fff94 ;
    memory[665] = 32'hbe1f566c ;
    memory[666] = 32'hbe258ba5 ;
    memory[667] = 32'h3de7321a ;
    memory[668] = 32'hbe066a4c ;
    memory[669] = 32'hbc960f95 ;
    memory[670] = 32'h3e0e2170 ;
    memory[671] = 32'h3e00ef5c ;
    memory[672] = 32'h3e0ed622 ;
    memory[673] = 32'hbdc29adc ;
    memory[674] = 32'h3cf18656 ;
    memory[675] = 32'h3da45bed ;
    memory[676] = 32'hbd373177 ;
    memory[677] = 32'hbd64223d ;
    memory[678] = 32'hbde7eaba ;
    memory[679] = 32'hbd40c530 ;
    memory[680] = 32'hbd525d3e ;
    memory[681] = 32'h3c8846b8 ;
    memory[682] = 32'hbda06cde ;
    memory[683] = 32'h3e1bb553 ;
    memory[684] = 32'h3d235a9a ;
    memory[685] = 32'h3dc7dd11 ;
    memory[686] = 32'hbc69b6c8 ;
    memory[687] = 32'hbd167331 ;
    memory[688] = 32'hbdfc131d ;
    memory[689] = 32'hbd86e9ea ;
    memory[690] = 32'hbd341ea7 ;
    memory[691] = 32'hbdd10034 ;
    memory[692] = 32'hbd546a4e ;
    memory[693] = 32'h3e08c72a ;
    memory[694] = 32'hbdb98b7a ;
    memory[695] = 32'h3e04d119 ;
    memory[696] = 32'hbd33448b ;
    memory[697] = 32'hbe13b508 ;
    memory[698] = 32'hbde7b206 ;
    memory[699] = 32'hbe020e9b ;
    memory[700] = 32'hbd9f9104 ;
    memory[701] = 32'hbd941b46 ;
    memory[702] = 32'h3e1045c8 ;
    memory[703] = 32'hbd9d9b7a ;
    memory[704] = 32'h3dd541ee ;
    memory[705] = 32'hbc370cf7 ;
    memory[706] = 32'h3d36ebd5 ;
    memory[707] = 32'hbd24da95 ;
    memory[708] = 32'hbd7cb973 ;
    memory[709] = 32'hbced1729 ;
    memory[710] = 32'h3d9a557a ;
    memory[711] = 32'h3d8efe57 ;
    memory[712] = 32'h3c43e5c9 ;
    memory[713] = 32'h3dafcd21 ;
    memory[714] = 32'h3e29881d ;
    memory[715] = 32'hbdf23fe6 ;
    memory[716] = 32'h3a625448 ;
    memory[717] = 32'h3e18c5b0 ;
    memory[718] = 32'h3da73433 ;
    memory[719] = 32'hbe14d104 ;
    memory[720] = 32'h3dadfc9f ;
    memory[721] = 32'hbd7e4cc3 ;
    memory[722] = 32'hbc7fe0cd ;
    memory[723] = 32'h3d556eb1 ;
    memory[724] = 32'hbd819cd9 ;
    memory[725] = 32'h3ca6c0b8 ;
    memory[726] = 32'h3ce67882 ;
    memory[727] = 32'hbe08bfe7 ;
    memory[728] = 32'h3d9e5bdb ;
    memory[729] = 32'h3dbdd3b3 ;
    memory[730] = 32'h3c36ccdd ;
    memory[731] = 32'h3dddadb8 ;
    memory[732] = 32'hbdad0423 ;
    memory[733] = 32'hbe0e2d03 ;
    memory[734] = 32'hbe358e66 ;
    memory[735] = 32'hbe0a9114 ;
    memory[736] = 32'h3ddf9f5e ;
    memory[737] = 32'hbdba2ce0 ;
    memory[738] = 32'h3d74da1e ;
    memory[739] = 32'hbd6aa29e ;
    memory[740] = 32'h3e040391 ;
    memory[741] = 32'hbd885375 ;
    memory[742] = 32'h3c618546 ;
    memory[743] = 32'hbca34f02 ;
    memory[744] = 32'h3e0904d7 ;
    memory[745] = 32'hbe02df99 ;
    memory[746] = 32'hbc2d4911 ;
    memory[747] = 32'h3e253842 ;
    memory[748] = 32'hbe16b7e5 ;
    memory[749] = 32'hbd12301e ;
    memory[750] = 32'h3e09aea7 ;
    memory[751] = 32'h3d453a56 ;
    memory[752] = 32'h3dda6ce1 ;
    memory[753] = 32'h3e074c46 ;
    memory[754] = 32'h3c8c48dd ;
    memory[755] = 32'hbbdcf65e ;
    memory[756] = 32'hbde8cbc7 ;
    memory[757] = 32'hbc51b88c ;
    memory[758] = 32'h3e3f688b ;
    memory[759] = 32'hbe204223 ;
    memory[760] = 32'hbde322ad ;
    memory[761] = 32'h3e21eb89 ;
    memory[762] = 32'hbe1d5e99 ;
    memory[763] = 32'hbd075d88 ;
    memory[764] = 32'h3d0e8571 ;
    memory[765] = 32'hbe49cd09 ;
    memory[766] = 32'hbc28a1ab ;
    memory[767] = 32'hbe187394 ;
    memory[768] = 32'h3d84dc9f ;
    memory[769] = 32'h3d10cd91 ;
    memory[770] = 32'hbe1ba613 ;
    memory[771] = 32'hbe274813 ;
    memory[772] = 32'hbe3e7c18 ;
    memory[773] = 32'h3e214454 ;
    memory[774] = 32'hbe0e3e13 ;
    memory[775] = 32'h3d93d33b ;
    memory[776] = 32'h3df9dd33 ;
    memory[777] = 32'h3cd1c2ce ;
    memory[778] = 32'hbb39de1b ;
    memory[779] = 32'h3d34c82f ;
    memory[780] = 32'h3df975b6 ;
    memory[781] = 32'hbe34af41 ;
    memory[782] = 32'h3e0c604b ;
    memory[783] = 32'h3e063d6e ;
    memory[784] = 32'hbd85af14 ;
    memory[785] = 32'hbcea3cef ;
    memory[786] = 32'h3d95821d ;
    memory[787] = 32'hbe1de9de ;
    memory[788] = 32'h3e017ce5 ;
    memory[789] = 32'hbe1b304d ;
    memory[790] = 32'h3d72cad4 ;
    memory[791] = 32'h3af72a57 ;
    memory[792] = 32'hbdf80a9a ;
    memory[793] = 32'h3e0ac740 ;
    memory[794] = 32'h3e235d70 ;
    memory[795] = 32'hbe0bc36c ;
    memory[796] = 32'hbdfbbd56 ;
    memory[797] = 32'h3a8e6991 ;
    memory[798] = 32'hbe265f0a ;
    memory[799] = 32'h3d612ce2 ;
    memory[800] = 32'hbd96bb15 ;
    memory[801] = 32'h3df9b700 ;
    memory[802] = 32'hbdb823d2 ;
    memory[803] = 32'h3b4d224a ;
    memory[804] = 32'hbdc5c94b ;
    memory[805] = 32'h3cb21354 ;
    memory[806] = 32'h3df49fe6 ;
    memory[807] = 32'h3d659599 ;
    memory[808] = 32'h3e2e0f0c ;
    memory[809] = 32'hbdab9c56 ;
    memory[810] = 32'hbe2b3655 ;
    memory[811] = 32'hbbc8c377 ;
    memory[812] = 32'h3e36fcf2 ;
    memory[813] = 32'h3da79eee ;
    memory[814] = 32'h3d3803d1 ;
    memory[815] = 32'h3dcc587a ;
    memory[816] = 32'h3d916a0a ;
    memory[817] = 32'h3e2ffaee ;
    memory[818] = 32'h3e0a4aaf ;
    memory[819] = 32'hbe298307 ;
    memory[820] = 32'hbccf72d8 ;
    memory[821] = 32'hbccfbefb ;
    memory[822] = 32'hbda016b8 ;
    memory[823] = 32'h3db9ed8c ;
    memory[824] = 32'hbdad0d56 ;
    memory[825] = 32'hbe07d2e3 ;
    memory[826] = 32'hbd56a391 ;
    memory[827] = 32'hbe150ce3 ;
    memory[828] = 32'hbdc405f2 ;
    memory[829] = 32'hbd9dc9b0 ;
    memory[830] = 32'hbe466251 ;
    memory[831] = 32'hbd12d5e1 ;
    memory[832] = 32'hbd4ddfc9 ;
    memory[833] = 32'hbe0677cd ;
    memory[834] = 32'h3d01e397 ;
    memory[835] = 32'h3c70b27e ;
    memory[836] = 32'h3e23624b ;
    memory[837] = 32'h3cc50879 ;
    memory[838] = 32'h3e113997 ;
    memory[839] = 32'h3e14e112 ;
    memory[840] = 32'h3cd3a409 ;
    memory[841] = 32'hbe32a6d5 ;
    memory[842] = 32'h3cbb24a4 ;
    memory[843] = 32'hbbdbe1df ;
    memory[844] = 32'h3e2fd1b5 ;
    memory[845] = 32'h3e09ac98 ;
    memory[846] = 32'hbdea6835 ;
    memory[847] = 32'h3dbcd08c ;
    memory[848] = 32'hbde1aef7 ;
    memory[849] = 32'h3e2c1375 ;
    memory[850] = 32'h3de02235 ;
    memory[851] = 32'hba098987 ;
    memory[852] = 32'h3d969263 ;
    memory[853] = 32'hbbae997d ;
    memory[854] = 32'h3df89042 ;
    memory[855] = 32'h3e05b4bf ;
    memory[856] = 32'hbe403143 ;
    memory[857] = 32'hbdbb7abc ;
    memory[858] = 32'h3d4580ea ;
    memory[859] = 32'h3d38546c ;
    memory[860] = 32'h3db658b4 ;
    memory[861] = 32'hbe22fc06 ;
    memory[862] = 32'hbd1daa7e ;
    memory[863] = 32'h3dc0719c ;
    memory[864] = 32'hbe1dca84 ;
    memory[865] = 32'hbc9061bb ;
    memory[866] = 32'h3e2c7daf ;
    memory[867] = 32'hbd42eaa7 ;
    memory[868] = 32'hbdb314f4 ;
    memory[869] = 32'h3d330c77 ;
    memory[870] = 32'h3d6b92c5 ;
    memory[871] = 32'h3d365f4a ;
    memory[872] = 32'h3d5f57c9 ;
    memory[873] = 32'hbe154be5 ;
    memory[874] = 32'h3de8340e ;
    memory[875] = 32'h3db2a5a0 ;
    memory[876] = 32'hbda0b468 ;
    memory[877] = 32'hbd0e8d47 ;
    memory[878] = 32'h3e19f085 ;
    memory[879] = 32'hbdbbc6aa ;
    memory[880] = 32'hbe04f3fa ;
    memory[881] = 32'hbde23d55 ;
    memory[882] = 32'hbd991c63 ;
    memory[883] = 32'hbdffe811 ;
    memory[884] = 32'hbd8d69b7 ;
    memory[885] = 32'hbdefa37e ;
    memory[886] = 32'h3d10cd1a ;
    memory[887] = 32'hba03fcf2 ;
    memory[888] = 32'h3c8feb9d ;
    memory[889] = 32'hbe2693d3 ;
    memory[890] = 32'h3d0bbbe0 ;
    memory[891] = 32'h3cac6c6f ;
    memory[892] = 32'hbdc62736 ;
    memory[893] = 32'hbe1ebe50 ;
    memory[894] = 32'hbd77e56c ;
    memory[895] = 32'h3e19ba5d ;
    memory[896] = 32'hbdcd12c0 ;
    memory[897] = 32'hbd728353 ;
    memory[898] = 32'h3e3ea6d1 ;
    memory[899] = 32'hbe1f3cfc ;
    memory[900] = 32'h3db81219 ;
    memory[901] = 32'hbe1f6376 ;
    memory[902] = 32'hbdaee23f ;
    memory[903] = 32'h3d8a8529 ;
    memory[904] = 32'hbdd40859 ;
    memory[905] = 32'h3c00325c ;
    memory[906] = 32'h3e1521b4 ;
    memory[907] = 32'hbe26af78 ;
    memory[908] = 32'h3dbea753 ;
    memory[909] = 32'hbd422967 ;
    memory[910] = 32'hbd3e9d7d ;
    memory[911] = 32'h3df39fd5 ;
    memory[912] = 32'hbdd72ec1 ;
    memory[913] = 32'hbd988321 ;
    memory[914] = 32'hbe112410 ;
    memory[915] = 32'hbd824909 ;
    memory[916] = 32'hbc465ef9 ;
    memory[917] = 32'h3c339911 ;
    memory[918] = 32'hbd852d70 ;
    memory[919] = 32'h3d9bb43b ;
    memory[920] = 32'hbe0c68d7 ;
    memory[921] = 32'hbbbdeb5e ;
    memory[922] = 32'h3d99b9a8 ;
    memory[923] = 32'h3e42c8fb ;
    memory[924] = 32'hbda8b932 ;
    memory[925] = 32'hbe164e54 ;
    memory[926] = 32'h3e1beb78 ;
    memory[927] = 32'h3dcca7f2 ;
    memory[928] = 32'hbde99920 ;
    memory[929] = 32'hbd86787e ;
    memory[930] = 32'hbdfb0db7 ;
    memory[931] = 32'h3cb970be ;
    memory[932] = 32'h3df25c3b ;
    memory[933] = 32'h3e14c59f ;
    memory[934] = 32'hbde146c3 ;
    memory[935] = 32'hbd086755 ;
    memory[936] = 32'hbd9814a5 ;
    memory[937] = 32'hbc1fbcb8 ;
    memory[938] = 32'h3d3d32f2 ;
    memory[939] = 32'h3d5ae6ee ;
    memory[940] = 32'h3e23b863 ;
    memory[941] = 32'hbddcbbcb ;
    memory[942] = 32'h3db0702c ;
    memory[943] = 32'hbdc4eada ;
    memory[944] = 32'hbd5ef147 ;
    memory[945] = 32'hbc163a94 ;
    memory[946] = 32'h3e2c9bb4 ;
    memory[947] = 32'hbd57d09e ;
    memory[948] = 32'hbd555884 ;
    memory[949] = 32'h3e1a6d2a ;
    memory[950] = 32'h3e2c64e1 ;
    memory[951] = 32'hbe1040d7 ;
    memory[952] = 32'h3e04fa3d ;
    memory[953] = 32'h3e11a685 ;
    memory[954] = 32'hbdbb7f43 ;
    memory[955] = 32'h3e1e7227 ;
    memory[956] = 32'hbe245009 ;
    memory[957] = 32'h3dd80c50 ;
    memory[958] = 32'hbe39dec0 ;
    memory[959] = 32'hbe2695e0 ;
    memory[960] = 32'hbe0003ce ;
    memory[961] = 32'hbdcdd067 ;
    memory[962] = 32'hbdcb4131 ;
    memory[963] = 32'hbdaf2e24 ;
    memory[964] = 32'h3e454344 ;
    memory[965] = 32'h3d99e6f5 ;
    memory[966] = 32'h3e09a786 ;
    memory[967] = 32'h3d5f6e6b ;
    memory[968] = 32'h3d237696 ;
    memory[969] = 32'h3e0de141 ;
    memory[970] = 32'h3da0862f ;
    memory[971] = 32'h3d2fe265 ;
    memory[972] = 32'h3df93b4b ;
    memory[973] = 32'hbd1e561b ;
    memory[974] = 32'hbd5109e2 ;
    memory[975] = 32'h3d4fdd6a ;
    memory[976] = 32'h3cc3e534 ;
    memory[977] = 32'hbdff30c6 ;
    memory[978] = 32'h3e114b84 ;
    memory[979] = 32'hbe18331b ;
    memory[980] = 32'h3d519aa0 ;
    memory[981] = 32'h3e292c1a ;
    memory[982] = 32'h3dc8e751 ;
    memory[983] = 32'h3c6089ed ;
    memory[984] = 32'h3c57f785 ;
    memory[985] = 32'hbd68d5b1 ;
    memory[986] = 32'hbd9f809c ;
    memory[987] = 32'h3da599c6 ;
    memory[988] = 32'hbdff4cb3 ;
    memory[989] = 32'h3dabf586 ;
    memory[990] = 32'h3d617d02 ;
    memory[991] = 32'hbd8480c3 ;
    memory[992] = 32'h3e052203 ;
    memory[993] = 32'hbdcd4037 ;
    memory[994] = 32'hbd9d4387 ;
    memory[995] = 32'h3bb83fac ;
    memory[996] = 32'h3cfabd15 ;
    memory[997] = 32'hbdcc8b5e ;
    memory[998] = 32'hbce2fc5d ;
    memory[999] = 32'h3d3ff59d ;
    memory[1000] = 32'hbe1ed55e ;
    memory[1001] = 32'hbd24a12c ;
    memory[1002] = 32'hbd7ca227 ;
    memory[1003] = 32'hbdc9c487 ;
    memory[1004] = 32'hbd9af865 ;
    memory[1005] = 32'h3bd6554e ;
    memory[1006] = 32'hbd407dad ;
    memory[1007] = 32'hbe2b5dfd ;
    memory[1008] = 32'hbe423c19 ;
    memory[1009] = 32'hbe15eff9 ;
    memory[1010] = 32'h3daee945 ;
    memory[1011] = 32'h3cc6f640 ;
    memory[1012] = 32'hbce7e7ee ;
    memory[1013] = 32'h3ccc8747 ;
    memory[1014] = 32'h3dd5c5f0 ;
    memory[1015] = 32'hbe06258f ;
    memory[1016] = 32'hbe03cfa9 ;
    memory[1017] = 32'h3e1aef30 ;
    memory[1018] = 32'h3d238537 ;
    memory[1019] = 32'h3d9454e8 ;
    memory[1020] = 32'h3e0eeb1d ;
    memory[1021] = 32'hbe19506c ;
    memory[1022] = 32'h3d8e8252 ;
    memory[1023] = 32'hbcccc1da ;
    memory[1024] = 32'hbdf88bb0 ;
    memory[1025] = 32'hbe2d16ff ;
    memory[1026] = 32'hbe0f6550 ;
    memory[1027] = 32'h3e389992 ;
    memory[1028] = 32'hbe2c9ec9 ;
    memory[1029] = 32'h3d13a61b ;
    memory[1030] = 32'h3e193064 ;
    memory[1031] = 32'h3e3c5f08 ;
    memory[1032] = 32'h3e07f16b ;
    memory[1033] = 32'hbe01f4a8 ;
    memory[1034] = 32'h3e3b7fb0 ;
    memory[1035] = 32'hbdacf720 ;
    memory[1036] = 32'h3e187ee3 ;
    memory[1037] = 32'h3e03d6ba ;
    memory[1038] = 32'h3d8334c7 ;
    memory[1039] = 32'hbe0cd860 ;
    memory[1040] = 32'hbdf7d707 ;
    memory[1041] = 32'hbe3bcfe0 ;
    memory[1042] = 32'hbe1776bf ;
    memory[1043] = 32'h3d4e7633 ;
    memory[1044] = 32'h3dcb2076 ;
    memory[1045] = 32'h3d9932ea ;
    memory[1046] = 32'h3de184a4 ;
    memory[1047] = 32'hbdd96ada ;
    memory[1048] = 32'h3e344de1 ;
    memory[1049] = 32'h3da01c78 ;
    memory[1050] = 32'h3e41c6c1 ;
    memory[1051] = 32'hbcda3ba8 ;
    memory[1052] = 32'h3d1d015f ;
    memory[1053] = 32'hbda75ea0 ;
    memory[1054] = 32'h3dd69928 ;
    memory[1055] = 32'hbe107e80 ;
    memory[1056] = 32'h3b9a3307 ;
    memory[1057] = 32'h3dcb78be ;
    memory[1058] = 32'hbdc7a4e9 ;
    memory[1059] = 32'h3cd94ff4 ;
    memory[1060] = 32'hbd04996d ;
    memory[1061] = 32'h3dbc32a0 ;
    memory[1062] = 32'hbd6786c7 ;
    memory[1063] = 32'hbadf6c18 ;
    memory[1064] = 32'h3cdfa272 ;
    memory[1065] = 32'hbc977458 ;
    memory[1066] = 32'hbd225316 ;
    memory[1067] = 32'hbdf96004 ;
    memory[1068] = 32'h3c8a1f4a ;
    memory[1069] = 32'hbd77464f ;
    memory[1070] = 32'h3db439e4 ;
    memory[1071] = 32'h3d959628 ;
    memory[1072] = 32'hbe19117e ;
    memory[1073] = 32'hbbb23e21 ;
    memory[1074] = 32'h3e159b8c ;
    memory[1075] = 32'hbdb66c79 ;
    memory[1076] = 32'h3cd8fdc1 ;
    memory[1077] = 32'h3dd88e1b ;
    memory[1078] = 32'hbe33ecf8 ;
    memory[1079] = 32'h3c28d557 ;
    memory[1080] = 32'h3cff992f ;
    memory[1081] = 32'h3e150d55 ;
    memory[1082] = 32'hbdcceeec ;
    memory[1083] = 32'h3dc55ace ;
    memory[1084] = 32'h3d80f2bb ;
    memory[1085] = 32'h3dbf72ed ;
    memory[1086] = 32'hbd02568b ;
    memory[1087] = 32'hbe0a6c3e ;
    memory[1088] = 32'h3cab72e4 ;
    memory[1089] = 32'hbd4683fd ;
    memory[1090] = 32'hbcaa8656 ;
    memory[1091] = 32'h3dde6863 ;
    memory[1092] = 32'hbe16c0b3 ;
    memory[1093] = 32'hbdac8a97 ;
    memory[1094] = 32'h3dfb1a2a ;
    memory[1095] = 32'h3e22dcd8 ;
    memory[1096] = 32'h3e1b3aa8 ;
    memory[1097] = 32'h3d0d3c4b ;
    memory[1098] = 32'h3dca07a8 ;
    memory[1099] = 32'h3d5f7e97 ;
    memory[1100] = 32'h3e3a0afb ;
    memory[1101] = 32'h3d8271e4 ;
    memory[1102] = 32'hbe1209ea ;
    memory[1103] = 32'hbe072efc ;
    memory[1104] = 32'hbc1588d3 ;
    memory[1105] = 32'h3ddf4399 ;
    memory[1106] = 32'hbe024eda ;
    memory[1107] = 32'h3e1fd146 ;
    memory[1108] = 32'h3e01d65a ;
    memory[1109] = 32'hbe27b2f9 ;
    memory[1110] = 32'hbe28acf7 ;
    memory[1111] = 32'hbdf3b5a8 ;
    memory[1112] = 32'hbdef1bd0 ;
    memory[1113] = 32'h3d5b6cfa ;
    memory[1114] = 32'h3d4c7e5c ;
    memory[1115] = 32'h3dc3037e ;
    memory[1116] = 32'hbb230a0a ;
    memory[1117] = 32'hbe029344 ;
    memory[1118] = 32'h3d1c5149 ;
    memory[1119] = 32'hbe17f8f8 ;
    memory[1120] = 32'hbd229921 ;
    memory[1121] = 32'h3c9718ec ;
    memory[1122] = 32'hbd9e07b3 ;
    memory[1123] = 32'hbbb8adde ;
    memory[1124] = 32'h3cbeaae5 ;
    memory[1125] = 32'h3d88aff2 ;
    memory[1126] = 32'hba7723cd ;
    memory[1127] = 32'hbdb02717 ;
    memory[1128] = 32'h3d97ba8f ;
    memory[1129] = 32'hbdac6def ;
    memory[1130] = 32'h3c3bf39b ;
    memory[1131] = 32'h3e22d35b ;
    memory[1132] = 32'hbe209d13 ;
    memory[1133] = 32'h3ccd4b35 ;
    memory[1134] = 32'h3dde8fe2 ;
    memory[1135] = 32'h3dc390bb ;
    memory[1136] = 32'hbc2923e6 ;
    memory[1137] = 32'hbd8d0300 ;
    memory[1138] = 32'h3cefafb2 ;
    memory[1139] = 32'h3dd43e46 ;
    memory[1140] = 32'h3d33ef15 ;
    memory[1141] = 32'h3c06d23f ;
    memory[1142] = 32'hbdd816e4 ;
    memory[1143] = 32'hbd6b7ba4 ;
    memory[1144] = 32'h3d4521ba ;
    memory[1145] = 32'hbdcdf9e8 ;
    memory[1146] = 32'h3cda78dd ;
    memory[1147] = 32'h3cb0da64 ;
    memory[1148] = 32'h3def9c0a ;
    memory[1149] = 32'h3df59f0b ;
    memory[1150] = 32'h3e01bba0 ;
    memory[1151] = 32'h3cfc3075 ;
    memory[1152] = 32'hbda5c6d7 ;
    memory[1153] = 32'h3aac180a ;
    memory[1154] = 32'h3e2049b2 ;
    memory[1155] = 32'hbc9108ae ;
    memory[1156] = 32'hbce2e279 ;
    memory[1157] = 32'hbc4d2012 ;
    memory[1158] = 32'h3e1f0d58 ;
    memory[1159] = 32'h3dc66fa7 ;
    memory[1160] = 32'h3d8f0020 ;
    memory[1161] = 32'hbe1f116d ;
    memory[1162] = 32'hbe00dedd ;
    memory[1163] = 32'h3c62dcdf ;
    memory[1164] = 32'h3e0d61f8 ;
    memory[1165] = 32'h3dd19ce1 ;
    memory[1166] = 32'hbdb221ac ;
    memory[1167] = 32'h3df7cceb ;
    memory[1168] = 32'hbdc33b65 ;
    memory[1169] = 32'h3e040c0b ;
    memory[1170] = 32'hbdf87a4d ;
    memory[1171] = 32'h3e00d510 ;
    memory[1172] = 32'h3caf07cd ;
    memory[1173] = 32'h3d303444 ;
    memory[1174] = 32'h3e37c270 ;
    memory[1175] = 32'hbe1d5ce3 ;
    memory[1176] = 32'h3da33a7f ;
    memory[1177] = 32'hbcc0e7a3 ;
    memory[1178] = 32'hbe069919 ;
    memory[1179] = 32'hbd6388c9 ;
    memory[1180] = 32'hbc8ebdf8 ;
    memory[1181] = 32'h3e2da444 ;
    memory[1182] = 32'hbe376264 ;
    memory[1183] = 32'hbcddc426 ;
    memory[1184] = 32'h3e0e50b9 ;
    memory[1185] = 32'hbd2e961f ;
    memory[1186] = 32'h3cfda13e ;
    memory[1187] = 32'hbd6fce62 ;
    memory[1188] = 32'h3e161008 ;
    memory[1189] = 32'h3dfdafe2 ;
    memory[1190] = 32'h3d2bbe27 ;
    memory[1191] = 32'hbdb883c1 ;
    memory[1192] = 32'hbdabcf66 ;
    memory[1193] = 32'h3e25f82b ;
    memory[1194] = 32'hbd5170c4 ;
    memory[1195] = 32'h3c6b3a74 ;
    memory[1196] = 32'hbdc4141a ;
    memory[1197] = 32'h3c0d6e7b ;
    memory[1198] = 32'h3e1fe104 ;
    memory[1199] = 32'h3d4772eb ;
    memory[1200] = 32'hbcf9d526 ;
    memory[1201] = 32'hbe2e5c69 ;
    memory[1202] = 32'h3bca1864 ;
    memory[1203] = 32'hbb7a96cb ;
    memory[1204] = 32'hbe1a2deb ;
    memory[1205] = 32'hbe243551 ;
    memory[1206] = 32'h3e3bdad4 ;
    memory[1207] = 32'hba2d8803 ;
    memory[1208] = 32'hbcf5709a ;
    memory[1209] = 32'h3ce82f11 ;
    memory[1210] = 32'hbe54a67b ;
    memory[1211] = 32'h3df0ac67 ;
    memory[1212] = 32'h3df30bbe ;
    memory[1213] = 32'h3ce1d170 ;
    memory[1214] = 32'h3db15686 ;
    memory[1215] = 32'hbdafd7b0 ;
    memory[1216] = 32'hbe16de57 ;
    memory[1217] = 32'h3d8cd3cc ;
    memory[1218] = 32'hbde2d4fa ;
    memory[1219] = 32'hbdd07570 ;
    memory[1220] = 32'h3e03be81 ;
    memory[1221] = 32'hbe019f94 ;
    memory[1222] = 32'hbe2db512 ;
    memory[1223] = 32'h3d8d85f9 ;
    memory[1224] = 32'h3e009a5a ;
    memory[1225] = 32'hbe2838cf ;
    memory[1226] = 32'hbd46577e ;
    memory[1227] = 32'h3e22f1a6 ;
    memory[1228] = 32'h3d11ecda ;
    memory[1229] = 32'hbdc850d5 ;
    memory[1230] = 32'hbde11ce9 ;
    memory[1231] = 32'hbe0c3216 ;
    memory[1232] = 32'hbe12ea29 ;
    memory[1233] = 32'h3de2049b ;
    memory[1234] = 32'hbd2a29b6 ;
    memory[1235] = 32'h3e07c93d ;
    memory[1236] = 32'hbdc40253 ;
    memory[1237] = 32'hbe0deb51 ;
    memory[1238] = 32'h3d4919db ;
    memory[1239] = 32'h3dd236ee ;
    memory[1240] = 32'hbc2d312f ;
    memory[1241] = 32'h3d01e968 ;
    memory[1242] = 32'hbe0b29c5 ;
    memory[1243] = 32'hbd2c0299 ;
    memory[1244] = 32'hbe28843e ;
    memory[1245] = 32'h3d51f96e ;
    memory[1246] = 32'h3c3c5333 ;
    memory[1247] = 32'hbda73eb9 ;
    memory[1248] = 32'hbcfd4e31 ;
    memory[1249] = 32'hbe1a180c ;
    memory[1250] = 32'hbe1c476c ;
    memory[1251] = 32'h3db187c3 ;
    memory[1252] = 32'hbc28270b ;
    memory[1253] = 32'h3e3dc6c5 ;
    memory[1254] = 32'h3d86b0f2 ;
    memory[1255] = 32'hbdf83270 ;
    memory[1256] = 32'hbdd01618 ;
    memory[1257] = 32'h3e2259b6 ;
    memory[1258] = 32'hbe3b1a69 ;
    memory[1259] = 32'h3d2b9a3b ;
    memory[1260] = 32'hbcdb2c02 ;
    memory[1261] = 32'hbd90a692 ;
    memory[1262] = 32'h3dcad956 ;
    memory[1263] = 32'hbd81b179 ;
    memory[1264] = 32'hbdda2aa6 ;
    memory[1265] = 32'h3d712ef4 ;
    memory[1266] = 32'hbd6f31d4 ;
    memory[1267] = 32'hbc269a6d ;
    memory[1268] = 32'hbca7755c ;
    memory[1269] = 32'h3e1d4f7f ;
    memory[1270] = 32'hbc2a4d46 ;
    memory[1271] = 32'h3e0cc3dc ;
    memory[1272] = 32'hbc775d1d ;
    memory[1273] = 32'hbe2c3de6 ;
    memory[1274] = 32'hbe10f5d3 ;
    memory[1275] = 32'hbd5248f5 ;
    memory[1276] = 32'h3e2a0176 ;
    memory[1277] = 32'h3c0d5373 ;
    memory[1278] = 32'h3e1b661e ;
    memory[1279] = 32'hbd6efa3f ;
    memory[1280] = 32'h3e437a44 ;
    memory[1281] = 32'h3e32f58a ;
    memory[1282] = 32'hbe017fab ;
    memory[1283] = 32'hbe19178a ;
    memory[1284] = 32'hbd66471d ;
    memory[1285] = 32'hbcf166d0 ;
    memory[1286] = 32'hbc8e1072 ;
    memory[1287] = 32'h3e291692 ;
    memory[1288] = 32'h3db0eb34 ;
    memory[1289] = 32'hbd87114f ;
    memory[1290] = 32'hbcbf966f ;
    memory[1291] = 32'hbe225f5b ;
    memory[1292] = 32'hbcfbfd72 ;
    memory[1293] = 32'hbe32b7b4 ;
    memory[1294] = 32'h3d22322c ;
    memory[1295] = 32'h3d9f1cf5 ;
    memory[1296] = 32'hbe1da7ec ;
    memory[1297] = 32'hbdaccbd2 ;
    memory[1298] = 32'h3e1ee87c ;
    memory[1299] = 32'hbe02f3b0 ;
    memory[1300] = 32'h3d273a90 ;
    memory[1301] = 32'h3daece69 ;
    memory[1302] = 32'h3d9fa1b8 ;
    memory[1303] = 32'hbe2ffddb ;
    memory[1304] = 32'hbe1accb4 ;
    memory[1305] = 32'hbe1cef5a ;
    memory[1306] = 32'h3dd8db27 ;
    memory[1307] = 32'h3ce78ccd ;
    memory[1308] = 32'h3da77870 ;
    memory[1309] = 32'hbdc4c0a8 ;
    memory[1310] = 32'hbdbfa5f4 ;
    memory[1311] = 32'hbe0c672e ;
    memory[1312] = 32'hbdb3f839 ;
    memory[1313] = 32'h3df0b173 ;
    memory[1314] = 32'hbdd7105a ;
    memory[1315] = 32'hbd5d0cb0 ;
    memory[1316] = 32'hbe072d35 ;
    memory[1317] = 32'hbd7d6623 ;
    memory[1318] = 32'h3e1a170a ;
    memory[1319] = 32'hbc7f2955 ;
    memory[1320] = 32'hbe315894 ;
    memory[1321] = 32'hbd9e0c17 ;
    memory[1322] = 32'hbdf6814e ;
    memory[1323] = 32'hbe049cad ;
    memory[1324] = 32'h3cdf9baf ;
    memory[1325] = 32'hba4e2ab7 ;
    memory[1326] = 32'h3d93f0bc ;
    memory[1327] = 32'hbcf1d8f8 ;
    memory[1328] = 32'h3e227f4f ;
    memory[1329] = 32'hbbd29d54 ;
    memory[1330] = 32'hbe18504e ;
    memory[1331] = 32'h3d741483 ;
    memory[1332] = 32'h3d3d179b ;
    memory[1333] = 32'hbcc99154 ;
    memory[1334] = 32'hbd25243d ;
    memory[1335] = 32'h3e47fc46 ;
    memory[1336] = 32'h3e4ebaab ;
    memory[1337] = 32'h3d7adc98 ;
    memory[1338] = 32'h3d029fc7 ;
    memory[1339] = 32'h3d22dd52 ;
    memory[1340] = 32'hbe101e4d ;
    memory[1341] = 32'h3e057323 ;
    memory[1342] = 32'hbca86083 ;
    memory[1343] = 32'h3e000193 ;
    memory[1344] = 32'h3e2e3899 ;
    memory[1345] = 32'hbdd00a1d ;
    memory[1346] = 32'hbe3fd619 ;
    memory[1347] = 32'hbcf4b91c ;
    memory[1348] = 32'h3e22f55a ;
    memory[1349] = 32'h3d18eb78 ;
    memory[1350] = 32'hbe11000e ;
    memory[1351] = 32'hbd58cabf ;
    memory[1352] = 32'hbd0401cd ;
    memory[1353] = 32'h3b9b578d ;
    memory[1354] = 32'hbe1d0169 ;
    memory[1355] = 32'h3d41a4a3 ;
    memory[1356] = 32'hbe31c0d5 ;
    memory[1357] = 32'hbc85a129 ;
    memory[1358] = 32'h3d51ecf0 ;
    memory[1359] = 32'h3e14b678 ;
    memory[1360] = 32'h3d002366 ;
    memory[1361] = 32'h3e22f247 ;
    memory[1362] = 32'h3dc7422d ;
    memory[1363] = 32'h3c50cf1e ;
    memory[1364] = 32'hbdc45831 ;
    memory[1365] = 32'hbd277738 ;
    memory[1366] = 32'h3dad60f3 ;
    memory[1367] = 32'hbde657a8 ;
    memory[1368] = 32'hbe62c6ef ;
    memory[1369] = 32'hbc4298e0 ;
    memory[1370] = 32'hbdff5c78 ;
    memory[1371] = 32'h3df4761b ;
    memory[1372] = 32'h3dd532f3 ;
    memory[1373] = 32'hbd8f3a71 ;
    memory[1374] = 32'h3dba76b1 ;
    memory[1375] = 32'h3db3175f ;
    memory[1376] = 32'hbe08c19d ;
    memory[1377] = 32'h3d843ac9 ;
    memory[1378] = 32'h3db3e417 ;
    memory[1379] = 32'h3dbe6f14 ;
    memory[1380] = 32'h39b3138c ;
    memory[1381] = 32'h3dc6daaf ;
    memory[1382] = 32'hbe24ec30 ;
    memory[1383] = 32'hbdccdcbf ;
    memory[1384] = 32'h3de459ae ;
    memory[1385] = 32'hbbd59a97 ;
    memory[1386] = 32'h3e2994ba ;
    memory[1387] = 32'hbdcac64c ;
    memory[1388] = 32'h3e12e4ab ;
    memory[1389] = 32'hbd3ed2f7 ;
    memory[1390] = 32'h3df6c334 ;
    memory[1391] = 32'h3e1b19bd ;
    memory[1392] = 32'h3d86b21c ;
    memory[1393] = 32'hbe32ad67 ;
    memory[1394] = 32'h3d04afc9 ;
    memory[1395] = 32'h3df0c8c8 ;
    memory[1396] = 32'h3d02e1a3 ;
    memory[1397] = 32'h3db05337 ;
    memory[1398] = 32'h3d8844c6 ;
    memory[1399] = 32'h3cadbfae ;
    memory[1400] = 32'hbdf38732 ;
    memory[1401] = 32'h3e01edd6 ;
    memory[1402] = 32'h3e6af945 ;
    memory[1403] = 32'hbdf3902f ;
    memory[1404] = 32'hbe0e2845 ;
    memory[1405] = 32'hbcf7942e ;
    memory[1406] = 32'hbc602015 ;
    memory[1407] = 32'hbdd2f49d ;
    memory[1408] = 32'h3d9fd0b5 ;
    memory[1409] = 32'h3d60e431 ;
    memory[1410] = 32'h3de37522 ;
    memory[1411] = 32'h3c31939e ;
    memory[1412] = 32'h3c315949 ;
    memory[1413] = 32'hbd83d735 ;
    memory[1414] = 32'h3d492d91 ;
    memory[1415] = 32'h3d96d526 ;
    memory[1416] = 32'hbcef20e1 ;
    memory[1417] = 32'hbdb5e94f ;
    memory[1418] = 32'hbd4ce495 ;
    memory[1419] = 32'h3de6c921 ;
    memory[1420] = 32'h3ddfc632 ;
    memory[1421] = 32'hbd927da4 ;
    memory[1422] = 32'hbe370bd6 ;
    memory[1423] = 32'hbc99737d ;
    memory[1424] = 32'h3aea5b71 ;
    memory[1425] = 32'h3e007a56 ;
    memory[1426] = 32'h3d04ad52 ;
    memory[1427] = 32'hbda3169f ;
    memory[1428] = 32'h3d40c529 ;
    memory[1429] = 32'hbc984712 ;
    memory[1430] = 32'hbc74284a ;
    memory[1431] = 32'h3db2e818 ;
    memory[1432] = 32'hbdb68ee9 ;
    memory[1433] = 32'h3d2ac132 ;
    memory[1434] = 32'hbdad928b ;
    memory[1435] = 32'h3dd9b338 ;
    memory[1436] = 32'h3e4842f4 ;
    memory[1437] = 32'h3dedb9ea ;
    memory[1438] = 32'hbbd44a4c ;
    memory[1439] = 32'h3d4e5af3 ;
    memory[1440] = 32'h3d9d3fa6 ;
    memory[1441] = 32'hbcaa4c7d ;
    memory[1442] = 32'hbbd49341 ;
    memory[1443] = 32'hbd91ee3f ;
    memory[1444] = 32'hbcc344ba ;
    memory[1445] = 32'hbe13a616 ;
    memory[1446] = 32'hbd7128be ;
    memory[1447] = 32'h3e26e697 ;
    memory[1448] = 32'h3db77ac1 ;
    memory[1449] = 32'hbe1fbd2f ;
    memory[1450] = 32'h3e11279f ;
    memory[1451] = 32'h3da178ab ;
    memory[1452] = 32'hbe0caf18 ;
    memory[1453] = 32'hbd950032 ;
    memory[1454] = 32'hbd926892 ;
    memory[1455] = 32'h3d7f71f3 ;
    memory[1456] = 32'h3de216ab ;
    memory[1457] = 32'hb87e71a4 ;
    memory[1458] = 32'h3d2caf32 ;
    memory[1459] = 32'hbc95dd61 ;
    memory[1460] = 32'h3c90a50c ;
    memory[1461] = 32'h3e23782c ;
    memory[1462] = 32'h3c0384cc ;
    memory[1463] = 32'h3c2c90e5 ;
    memory[1464] = 32'h3e2aff99 ;
    memory[1465] = 32'hbde588b5 ;
    memory[1466] = 32'hbd69052f ;
    memory[1467] = 32'h3d553044 ;
    memory[1468] = 32'hbd8faeb3 ;
    memory[1469] = 32'hbe241f38 ;
    memory[1470] = 32'hbe0961b2 ;
    memory[1471] = 32'h3de66da9 ;
    memory[1472] = 32'h3c9dc73f ;
    memory[1473] = 32'h3dfa9060 ;
    memory[1474] = 32'hbdc57de9 ;
    memory[1475] = 32'hbdfb80e8 ;
    memory[1476] = 32'hbe24f4e8 ;
    memory[1477] = 32'hbe1463a1 ;
    memory[1478] = 32'hbcfb9e46 ;
    memory[1479] = 32'h3e3becd2 ;
    memory[1480] = 32'h3cddc400 ;
    memory[1481] = 32'h3d2a3726 ;
    memory[1482] = 32'h3d81f9f9 ;
    memory[1483] = 32'h3dc649bd ;
    memory[1484] = 32'h3da021ff ;
    memory[1485] = 32'hbe0c0df2 ;
    memory[1486] = 32'hbd17d10a ;
    memory[1487] = 32'h3e0ae2e8 ;
    memory[1488] = 32'h3e143f22 ;
    memory[1489] = 32'h3daffe16 ;
    memory[1490] = 32'h3d40b343 ;
    memory[1491] = 32'h3d7453a7 ;
    memory[1492] = 32'hbdfbbf9b ;
    memory[1493] = 32'hbc91bb66 ;
    memory[1494] = 32'hbd9a55b5 ;
    memory[1495] = 32'h3db36271 ;
    memory[1496] = 32'h3e165056 ;
    memory[1497] = 32'hbded76bf ;
    memory[1498] = 32'h3dcbcb7d ;
    memory[1499] = 32'h3e3d5762 ;
    memory[1500] = 32'h3dad1429 ;
    memory[1501] = 32'hbdb47eb6 ;
    memory[1502] = 32'h3c9b0bc2 ;
    memory[1503] = 32'h3e3460ed ;
    memory[1504] = 32'hb94c4642 ;
    memory[1505] = 32'h3cd1869a ;
    memory[1506] = 32'h3da0e950 ;
    memory[1507] = 32'h3dfbaafc ;
    memory[1508] = 32'hbdc2d531 ;
    memory[1509] = 32'h3d1a102d ;
    memory[1510] = 32'h3cda429a ;
    memory[1511] = 32'h3cbd6b17 ;
    memory[1512] = 32'hbcd4e7e1 ;
    memory[1513] = 32'h3debb9d1 ;
    memory[1514] = 32'h3dcc5df2 ;
    memory[1515] = 32'hbe0850cb ;
    memory[1516] = 32'hbd9a3b2f ;
    memory[1517] = 32'hbd95cadb ;
    memory[1518] = 32'hbe0c28c4 ;
    memory[1519] = 32'h3db129fd ;
    memory[1520] = 32'h3dbb6b0d ;
    memory[1521] = 32'hbdf7aafb ;
    memory[1522] = 32'h3db5005d ;
    memory[1523] = 32'h3e35245f ;
    memory[1524] = 32'h3e065a5f ;
    memory[1525] = 32'hbdc026c8 ;
    memory[1526] = 32'h39a0fe93 ;
    memory[1527] = 32'h3d75b9be ;
    memory[1528] = 32'h3da4a2e5 ;
    memory[1529] = 32'h3d2aa03e ;
    memory[1530] = 32'hbe27f682 ;
    memory[1531] = 32'h3d38a599 ;
    memory[1532] = 32'h3ce28941 ;
    memory[1533] = 32'h3dcd81f6 ;
    memory[1534] = 32'hbd9de864 ;
    memory[1535] = 32'h3dafb0e1 ;
    memory[1536] = 32'h3e2be798 ;
    memory[1537] = 32'hbd4a47de ;
    memory[1538] = 32'h3c998482 ;
    memory[1539] = 32'h3d85a6ad ;
    memory[1540] = 32'hbe2df87a ;
    memory[1541] = 32'hbc29d23d ;
    memory[1542] = 32'h3dd0430a ;
    memory[1543] = 32'h3d11b7dd ;
    memory[1544] = 32'h3dc5215a ;
    memory[1545] = 32'h3e22deae ;
    memory[1546] = 32'h3e0a2f03 ;
    memory[1547] = 32'hbdbe5a8e ;
    memory[1548] = 32'h3df8c84c ;
    memory[1549] = 32'hbe1861b3 ;
    memory[1550] = 32'hbde83eb0 ;
    memory[1551] = 32'hbd371967 ;
    memory[1552] = 32'hbba3a83f ;
    memory[1553] = 32'h3e1096f4 ;
    memory[1554] = 32'h3e20f152 ;
    memory[1555] = 32'hbdd0ac92 ;
    memory[1556] = 32'hbdae69fc ;
    memory[1557] = 32'h3ce79dbc ;
    memory[1558] = 32'hbadfc105 ;
    memory[1559] = 32'h3d7cb40e ;
    memory[1560] = 32'hbdadf6fb ;
    memory[1561] = 32'hbdf98ffe ;
    memory[1562] = 32'hbcb17c58 ;
    memory[1563] = 32'h3e34484e ;
    memory[1564] = 32'h3d464e00 ;
    memory[1565] = 32'hbdb40cbd ;
    memory[1566] = 32'h3d6104d3 ;
    memory[1567] = 32'hbdd3a44b ;
    memory[1568] = 32'hbde8680c ;
    memory[1569] = 32'h3e1ed6f5 ;
    memory[1570] = 32'hb98f8614 ;
    memory[1571] = 32'h3d5b5070 ;
    memory[1572] = 32'h3d9bf08c ;
    memory[1573] = 32'hbd8b8e96 ;
    memory[1574] = 32'hbda298d4 ;
    memory[1575] = 32'hbd9eccb7 ;
    memory[1576] = 32'hbe1494a6 ;
    memory[1577] = 32'hbc8d4364 ;
    memory[1578] = 32'hbb52af24 ;
    memory[1579] = 32'hbdea31a6 ;
    memory[1580] = 32'h3e09938e ;
    memory[1581] = 32'hbe2cb0e4 ;
    memory[1582] = 32'h3e0bc04d ;
    memory[1583] = 32'h3e136dfe ;
    memory[1584] = 32'hbe29c847 ;
    memory[1585] = 32'hbe2a82f4 ;
    memory[1586] = 32'h3e297e76 ;
    memory[1587] = 32'hbcdce46e ;
    memory[1588] = 32'h3cb7f2d9 ;
    memory[1589] = 32'h3b4204a6 ;
    memory[1590] = 32'h3e131b4f ;
    memory[1591] = 32'hbd54c597 ;
    memory[1592] = 32'h3b6ec38b ;
    memory[1593] = 32'hbdcd5c56 ;
    memory[1594] = 32'h3df103de ;
    memory[1595] = 32'hbd9a5a2b ;
    memory[1596] = 32'h3dc3398a ;
    memory[1597] = 32'hbde35fa9 ;
    memory[1598] = 32'h3e0bb958 ;
    memory[1599] = 32'hbda18111 ;
    memory[1600] = 32'hbe12aa06 ;
    memory[1601] = 32'hbe1d4769 ;
    memory[1602] = 32'hbdd6c6ea ;
    memory[1603] = 32'hbc7ea65b ;
    memory[1604] = 32'hbe0ef28b ;
    memory[1605] = 32'h3e044487 ;
    memory[1606] = 32'h3d949757 ;
    memory[1607] = 32'h3e1976f6 ;
    memory[1608] = 32'hbda9ac8d ;
    memory[1609] = 32'h3e0dcbe2 ;
    memory[1610] = 32'h3e21e083 ;
    memory[1611] = 32'hbd627b34 ;
    memory[1612] = 32'hbd262b20 ;
    memory[1613] = 32'h3e14b6dd ;
    memory[1614] = 32'h3e4099b0 ;
    memory[1615] = 32'hbe14d1ea ;
    memory[1616] = 32'h3e1fe53f ;
    memory[1617] = 32'h3de2f07c ;
    memory[1618] = 32'h3e2d777f ;
    memory[1619] = 32'hbd5fcfda ;
    memory[1620] = 32'h3d4876c7 ;
    memory[1621] = 32'hbd814114 ;
    memory[1622] = 32'hbe2a83ba ;
    memory[1623] = 32'h3e32a4dd ;
    memory[1624] = 32'h3e34bcc3 ;
    memory[1625] = 32'hbe1def6a ;
    memory[1626] = 32'hbe018e20 ;
    memory[1627] = 32'h3d4f693e ;
    memory[1628] = 32'h3e142f76 ;
    memory[1629] = 32'hbd75d397 ;
    memory[1630] = 32'hbe06865d ;
    memory[1631] = 32'h3c161f6d ;
    memory[1632] = 32'h3d9c580d ;
    memory[1633] = 32'h3d3ffb93 ;
    memory[1634] = 32'h3e1a8bb6 ;
    memory[1635] = 32'h3e37cfe1 ;
    memory[1636] = 32'h3cedefa6 ;
    memory[1637] = 32'h3d8d4d4c ;
    memory[1638] = 32'hbd424827 ;
    memory[1639] = 32'h3d88c39f ;
    memory[1640] = 32'hbdb449fa ;
    memory[1641] = 32'h3dd1ba21 ;
    memory[1642] = 32'h3d068091 ;
    memory[1643] = 32'hbccd5911 ;
    memory[1644] = 32'h3d0e6c59 ;
    memory[1645] = 32'hbdcaa01a ;
    memory[1646] = 32'h3d7b6a57 ;
    memory[1647] = 32'hbd3d1e34 ;
    memory[1648] = 32'h3d6ea6ef ;
    memory[1649] = 32'hbd753a1d ;
    memory[1650] = 32'h3d3e3ce0 ;
    memory[1651] = 32'h3e0c1648 ;
    memory[1652] = 32'hbdc6c478 ;
    memory[1653] = 32'hbdf10d9c ;
    memory[1654] = 32'hbce23044 ;
    memory[1655] = 32'hbe28e2ba ;
    memory[1656] = 32'h3d3881fa ;
    memory[1657] = 32'h3c0247b0 ;
    memory[1658] = 32'hbda8d5a0 ;
    memory[1659] = 32'h3d35b5b4 ;
    memory[1660] = 32'hbd806da2 ;
    memory[1661] = 32'hbcc86753 ;
    memory[1662] = 32'h3e052dd5 ;
    memory[1663] = 32'hbd6f7791 ;
    memory[1664] = 32'hbdfb8802 ;
    memory[1665] = 32'hbe22ede9 ;
    memory[1666] = 32'h3d9fc973 ;
    memory[1667] = 32'h3d8a3a2b ;
    memory[1668] = 32'hbce6e2b3 ;
    memory[1669] = 32'hbe4247cb ;
    memory[1670] = 32'hbe2627d8 ;
    memory[1671] = 32'h3db844a5 ;
    memory[1672] = 32'hbdcab7eb ;
    memory[1673] = 32'h3dd406c6 ;
    memory[1674] = 32'h3ccf6478 ;
    memory[1675] = 32'hbd2b0586 ;
    memory[1676] = 32'hbe24534c ;
    memory[1677] = 32'h3e1f4448 ;
    memory[1678] = 32'hbc7a9a62 ;
    memory[1679] = 32'hbb0b5ed6 ;
    memory[1680] = 32'hbddffdb1 ;
    memory[1681] = 32'hbcafd236 ;
    memory[1682] = 32'hbcdd4378 ;
    memory[1683] = 32'h3e26663e ;
    memory[1684] = 32'h3dc3e050 ;
    memory[1685] = 32'hbdb0af4f ;
    memory[1686] = 32'h3d81f8c2 ;
    memory[1687] = 32'h3dd6d3f2 ;
    memory[1688] = 32'h3d0b9c1d ;
    memory[1689] = 32'hbd8f5f24 ;
    memory[1690] = 32'hbe01f79c ;
    memory[1691] = 32'hbe1d12ed ;
    memory[1692] = 32'hbd6e4e6d ;
    memory[1693] = 32'h3e17b084 ;
    memory[1694] = 32'hbd3878c9 ;
    memory[1695] = 32'hbe0d3f7d ;
    memory[1696] = 32'hbde6e743 ;
    memory[1697] = 32'hbc987038 ;
    memory[1698] = 32'hbd060d4a ;
    memory[1699] = 32'hbdb6fb72 ;
    memory[1700] = 32'h3d5b15df ;
    memory[1701] = 32'h3e21c775 ;
    memory[1702] = 32'h3bd9a4f8 ;
    memory[1703] = 32'h3d9d105c ;
    memory[1704] = 32'h3e30cd54 ;
    memory[1705] = 32'hbe128731 ;
    memory[1706] = 32'hbd3105b7 ;
    memory[1707] = 32'h3d72a218 ;
    memory[1708] = 32'h3e14dc27 ;
    memory[1709] = 32'h3dbb6940 ;
    memory[1710] = 32'hbc5248f8 ;
    memory[1711] = 32'hbdb12092 ;
    memory[1712] = 32'hbddfb46f ;
    memory[1713] = 32'hbd02aaf7 ;
    memory[1714] = 32'h3dbe37f2 ;
    memory[1715] = 32'hbda7b61a ;
    memory[1716] = 32'h3e21f442 ;
    memory[1717] = 32'h3d1dd38b ;
    memory[1718] = 32'h3de7f89d ;
    memory[1719] = 32'hbe2a7531 ;
    memory[1720] = 32'h3cdc383d ;
    memory[1721] = 32'h3d268810 ;
    memory[1722] = 32'hb9b0c7b1 ;
    memory[1723] = 32'hbd7e436a ;
    memory[1724] = 32'hbe33b1a4 ;
    memory[1725] = 32'h3dacf01a ;
    memory[1726] = 32'hbdb49315 ;
    memory[1727] = 32'hbe2861e4 ;
    memory[1728] = 32'h3de34574 ;
    memory[1729] = 32'h3e081fb5 ;
    memory[1730] = 32'hbdbdc1eb ;
    memory[1731] = 32'h3ccd07ac ;
    memory[1732] = 32'h3dfa1dfa ;
    memory[1733] = 32'hbcfebb42 ;
    memory[1734] = 32'h3c618c28 ;
    memory[1735] = 32'hbdd1694b ;
    memory[1736] = 32'hbd4bac2b ;
    memory[1737] = 32'h3e0a64f5 ;
    memory[1738] = 32'h3de163f1 ;
    memory[1739] = 32'hbe12c18a ;
    memory[1740] = 32'hbd978bf9 ;
    memory[1741] = 32'h3d853620 ;
    memory[1742] = 32'hbdcab197 ;
    memory[1743] = 32'hbe2212cb ;
    memory[1744] = 32'hbdbf879b ;
    memory[1745] = 32'h3dc5370f ;
    memory[1746] = 32'h3d34b797 ;
    memory[1747] = 32'hbdead1fc ;
    memory[1748] = 32'hbd4c0973 ;
    memory[1749] = 32'h3e0b07d9 ;
    memory[1750] = 32'hbd90f1de ;
    memory[1751] = 32'hbd90bfec ;
    memory[1752] = 32'h3cd954d4 ;
    memory[1753] = 32'hbc4a27ce ;
    memory[1754] = 32'hbe1183ef ;
    memory[1755] = 32'h3dd587ee ;
    memory[1756] = 32'hbd944cba ;
    memory[1757] = 32'h3e02d58f ;
    memory[1758] = 32'h3e1cfc10 ;
    memory[1759] = 32'h3de42e0d ;
    memory[1760] = 32'hbe1ccc13 ;
    memory[1761] = 32'hbbeb4cb2 ;
    memory[1762] = 32'h3dd3fc0b ;
    memory[1763] = 32'h3e3ee38a ;
    memory[1764] = 32'hbd43098a ;
    memory[1765] = 32'hbcccbe16 ;
    memory[1766] = 32'h3cb99d9d ;
    memory[1767] = 32'hbdd729a1 ;
    memory[1768] = 32'hbdef178f ;
    memory[1769] = 32'hbd811ae8 ;
    memory[1770] = 32'h3d10756d ;
    memory[1771] = 32'h3e150457 ;
    memory[1772] = 32'hbe694364 ;
    memory[1773] = 32'h3e2a180f ;
    memory[1774] = 32'hbdec4677 ;
    memory[1775] = 32'hbdba78d5 ;
    memory[1776] = 32'h3d1d00d2 ;
    memory[1777] = 32'h3d748248 ;
    memory[1778] = 32'h3e0b1625 ;
    memory[1779] = 32'h3e13069e ;
    memory[1780] = 32'hbde8b9bb ;
    memory[1781] = 32'h3e3aa6f8 ;
    memory[1782] = 32'hbd2836c9 ;
    memory[1783] = 32'h3d551497 ;
    memory[1784] = 32'h3e2edb9e ;
    memory[1785] = 32'hbc4cd0ad ;
    memory[1786] = 32'hbbec7bb3 ;
    memory[1787] = 32'hbc33f519 ;
    memory[1788] = 32'h3c96db0a ;
    memory[1789] = 32'hbe232d9e ;
    memory[1790] = 32'h3d8a833a ;
    memory[1791] = 32'hbd2ae8a9 ;
    memory[1792] = 32'hbda49743 ;
    memory[1793] = 32'h3d1f3087 ;
    memory[1794] = 32'hbd8c0b6d ;
    memory[1795] = 32'h3e13be9a ;
    memory[1796] = 32'h3d0f1ce8 ;
    memory[1797] = 32'h3e3b23a1 ;
    memory[1798] = 32'h3e1f3dac ;
    memory[1799] = 32'h3b74430d ;
    memory[1800] = 32'hbce6978d ;
    memory[1801] = 32'hbc8efca8 ;
    memory[1802] = 32'h3d885761 ;
    memory[1803] = 32'hbe12704f ;
    memory[1804] = 32'hbe07ee49 ;
    memory[1805] = 32'h3d99ef1d ;
    memory[1806] = 32'h3c91a155 ;
    memory[1807] = 32'h3e1d955c ;
    memory[1808] = 32'hbdd646c7 ;
    memory[1809] = 32'h3c73071f ;
    memory[1810] = 32'h3e5691bf ;
    memory[1811] = 32'h3dfb6b58 ;
    memory[1812] = 32'h3d3a0d91 ;
    memory[1813] = 32'hbe29a2d7 ;
    memory[1814] = 32'h3e3f5c13 ;
    memory[1815] = 32'hbd81e12b ;
    memory[1816] = 32'hbd7e6f67 ;
    memory[1817] = 32'hbd65c42a ;
    memory[1818] = 32'hbd841ac3 ;
    memory[1819] = 32'hbe06b014 ;
    memory[1820] = 32'h3c14d5dd ;
    memory[1821] = 32'h3e1fce51 ;
    memory[1822] = 32'hbd98cd96 ;
    memory[1823] = 32'hbd5247f0 ;
    memory[1824] = 32'hbe1c529c ;
    memory[1825] = 32'h3e140bc2 ;
    memory[1826] = 32'hbdf79be6 ;
    memory[1827] = 32'h3e2dd7d1 ;
    memory[1828] = 32'h3c769832 ;
    memory[1829] = 32'hbe06908b ;
    memory[1830] = 32'h3d51c73d ;
    memory[1831] = 32'hbd84496d ;
    memory[1832] = 32'hbdd95308 ;
    memory[1833] = 32'hbd635cc9 ;
    memory[1834] = 32'hbe03ed04 ;
    memory[1835] = 32'h3c8b44de ;
    memory[1836] = 32'hbd770ede ;
    memory[1837] = 32'hbdcfbdb4 ;
    memory[1838] = 32'h3da96035 ;
    memory[1839] = 32'hbdf8c3e5 ;
    memory[1840] = 32'hbd3c8f87 ;
    memory[1841] = 32'hbe19649a ;
    memory[1842] = 32'hbe2fcd10 ;
    memory[1843] = 32'hbde38c74 ;
    memory[1844] = 32'hbd8c5549 ;
    memory[1845] = 32'hbe0f7932 ;
    memory[1846] = 32'h3d270093 ;
    memory[1847] = 32'hbd811ac7 ;
    memory[1848] = 32'h3df5c2af ;
    memory[1849] = 32'h3e3e5940 ;
    memory[1850] = 32'h3dafad04 ;
    memory[1851] = 32'hbd23d730 ;
    memory[1852] = 32'h3e1bf8d5 ;
    memory[1853] = 32'hbdcd3224 ;
    memory[1854] = 32'hbe0439bf ;
    memory[1855] = 32'hbdba9206 ;
    memory[1856] = 32'hbdee0a04 ;
    memory[1857] = 32'h3dff446b ;
    memory[1858] = 32'h3cc11085 ;
    memory[1859] = 32'h3db16d3b ;
    memory[1860] = 32'h3d0089f0 ;
    memory[1861] = 32'hbe006e9d ;
    memory[1862] = 32'hbd7280d6 ;
    memory[1863] = 32'h3d7f356c ;
    memory[1864] = 32'hbe14281c ;
    memory[1865] = 32'h3d5ba286 ;
    memory[1866] = 32'h3d3716e7 ;
    memory[1867] = 32'h38411446 ;
    memory[1868] = 32'h3da6295d ;
    memory[1869] = 32'hbdc134c3 ;
    memory[1870] = 32'h3d700813 ;
    memory[1871] = 32'hbcbc9e25 ;
    memory[1872] = 32'hbd99b9bb ;
    memory[1873] = 32'hbe3c0bc6 ;
    memory[1874] = 32'hbdc9de32 ;
    memory[1875] = 32'h3e263a38 ;
    memory[1876] = 32'hbdf3f9f0 ;
    memory[1877] = 32'hbd8d20c2 ;
    memory[1878] = 32'hbe1adc01 ;
    memory[1879] = 32'h3e31c4b3 ;
    memory[1880] = 32'h3e361697 ;
    memory[1881] = 32'h3d07e298 ;
    memory[1882] = 32'hbc10c67f ;
    memory[1883] = 32'hbe301206 ;
    memory[1884] = 32'h3d9009bd ;
    memory[1885] = 32'hbd1c6b3c ;
    memory[1886] = 32'h3da5c7ad ;
    memory[1887] = 32'h3e1529e6 ;
    memory[1888] = 32'h3e156e2c ;
    memory[1889] = 32'hbe343390 ;
    memory[1890] = 32'h3e3c9307 ;
    memory[1891] = 32'hbdd5ea38 ;
    memory[1892] = 32'h3cfa8802 ;
    memory[1893] = 32'hbd46c1de ;
    memory[1894] = 32'h3e03d9de ;
    memory[1895] = 32'hbd38023a ;
    memory[1896] = 32'h3dd6daa9 ;
    memory[1897] = 32'hbcc7f093 ;
    memory[1898] = 32'hbd6c33df ;
    memory[1899] = 32'hbc856925 ;
    memory[1900] = 32'hbe102955 ;
    memory[1901] = 32'h3dbe8afe ;
    memory[1902] = 32'h3e53dec0 ;
    memory[1903] = 32'hbd627385 ;
    memory[1904] = 32'hbd1c9af8 ;
    memory[1905] = 32'hbdf88848 ;
    memory[1906] = 32'h3d9d0a11 ;
    memory[1907] = 32'hbbc2cf7c ;
    memory[1908] = 32'hbe242f34 ;
    memory[1909] = 32'h3dadff7f ;
    memory[1910] = 32'h3c41d848 ;
    memory[1911] = 32'h3e0efc6c ;
    memory[1912] = 32'hbd4e2b00 ;
    memory[1913] = 32'h3e15caa2 ;
    memory[1914] = 32'h3dc8e03d ;
    memory[1915] = 32'h3d0c12db ;
    memory[1916] = 32'h3e11b2cf ;
    memory[1917] = 32'hbe12d85a ;
    memory[1918] = 32'h3d0fe109 ;
    memory[1919] = 32'hbd55bb4b ;
    memory[1920] = 32'h3c1b47dc ;
    memory[1921] = 32'hbe237fe6 ;
    memory[1922] = 32'hbd169ee6 ;
    memory[1923] = 32'hbe1c2e8e ;
    memory[1924] = 32'hbdf7aff1 ;
    memory[1925] = 32'hbe50313e ;
    memory[1926] = 32'h3dd9d347 ;
    memory[1927] = 32'hbc3702be ;
    memory[1928] = 32'hbbca364e ;
    memory[1929] = 32'hbbf88f88 ;
    memory[1930] = 32'hbd353d17 ;
    memory[1931] = 32'h3d35fe7d ;
    memory[1932] = 32'hbc7e2b79 ;
    memory[1933] = 32'hbe2c3f00 ;
    memory[1934] = 32'h388f0da5 ;
    memory[1935] = 32'hbd022d95 ;
    memory[1936] = 32'h3d938792 ;
    memory[1937] = 32'hbe13b340 ;
    memory[1938] = 32'h3e198c27 ;
    memory[1939] = 32'h3d55c993 ;
    memory[1940] = 32'hbb03cd99 ;
    memory[1941] = 32'hbe01ab23 ;
    memory[1942] = 32'hbd57aad9 ;
    memory[1943] = 32'h3e26d334 ;
    memory[1944] = 32'h3de461d4 ;
    memory[1945] = 32'h3e430038 ;
    memory[1946] = 32'h3dd57492 ;
    memory[1947] = 32'h3e2d6799 ;
    memory[1948] = 32'h3ce08b01 ;
    memory[1949] = 32'hbd7711e5 ;
    memory[1950] = 32'h3d549ba6 ;
    memory[1951] = 32'h3e07cd66 ;
    memory[1952] = 32'h3ddb501b ;
    memory[1953] = 32'h3dd2e9a0 ;
    memory[1954] = 32'h3e161223 ;
    memory[1955] = 32'h3df51510 ;
    memory[1956] = 32'h3c2b07c8 ;
    memory[1957] = 32'h3e2d1871 ;
    memory[1958] = 32'h3d07498c ;
    memory[1959] = 32'h3da5a74f ;
    memory[1960] = 32'h3d09d5ca ;
    memory[1961] = 32'h3dc4557c ;
    memory[1962] = 32'h3e257422 ;
    memory[1963] = 32'h3c99e100 ;
    memory[1964] = 32'hbd4258f0 ;
    memory[1965] = 32'h3e2a357c ;
    memory[1966] = 32'h3d341225 ;
    memory[1967] = 32'h3decc9db ;
    memory[1968] = 32'h3c43cd49 ;
    memory[1969] = 32'hbcaebba5 ;
    memory[1970] = 32'hbe36c42a ;
    memory[1971] = 32'hbc993e66 ;
    memory[1972] = 32'h3db89068 ;
    memory[1973] = 32'h3c36317e ;
    memory[1974] = 32'h3d8d1360 ;
    memory[1975] = 32'hbe14c084 ;
    memory[1976] = 32'hbd21e206 ;
    memory[1977] = 32'hbd8ce80e ;
    memory[1978] = 32'hbde91c77 ;
    memory[1979] = 32'hbe183ebb ;
    memory[1980] = 32'hbe2f50e7 ;
    memory[1981] = 32'h3d6db6da ;
    memory[1982] = 32'hbd8a8270 ;
    memory[1983] = 32'h3dc7de89 ;
    memory[1984] = 32'h3e4b4ea7 ;
    memory[1985] = 32'h3c618eda ;
    memory[1986] = 32'hbe04b3c3 ;
    memory[1987] = 32'h3e197f7a ;
    memory[1988] = 32'h3ba018c1 ;
    memory[1989] = 32'h3d5740dc ;
    memory[1990] = 32'h3df37753 ;
    memory[1991] = 32'h3dbe8a82 ;
    memory[1992] = 32'h3e0e76eb ;
    memory[1993] = 32'hbdff9c77 ;
    memory[1994] = 32'h3e13029f ;
    memory[1995] = 32'h3e2208fe ;
    memory[1996] = 32'h3d13de02 ;
    memory[1997] = 32'hbd6377c3 ;
    memory[1998] = 32'hbe25178f ;
    memory[1999] = 32'hbe08e4ee ;
    memory[2000] = 32'h3dcf13a5 ;
    memory[2001] = 32'h3e27bd29 ;
    memory[2002] = 32'hbb5327c5 ;
    memory[2003] = 32'hbe252673 ;
    memory[2004] = 32'h3e39c8b0 ;
    memory[2005] = 32'h3d8f5528 ;
    memory[2006] = 32'hbdf7bc94 ;
    memory[2007] = 32'h3ce0692c ;
    memory[2008] = 32'h3d002fe0 ;
    memory[2009] = 32'h3cb5162c ;
    memory[2010] = 32'hbe29984c ;
    memory[2011] = 32'h3d73112c ;
    memory[2012] = 32'h3e1f7e71 ;
    memory[2013] = 32'hbe04c3aa ;
    memory[2014] = 32'h3dce4fee ;
    memory[2015] = 32'hbd24517a ;
    memory[2016] = 32'hbcb35607 ;
    memory[2017] = 32'hbd60f2db ;
    memory[2018] = 32'hbddcc4b9 ;
    memory[2019] = 32'hbe0ff400 ;
    memory[2020] = 32'hbe0b48a9 ;
    memory[2021] = 32'hbde63c47 ;
    memory[2022] = 32'hbbc4453b ;
    memory[2023] = 32'hbcf3cbd4 ;
    memory[2024] = 32'h3e08d08c ;
    memory[2025] = 32'h3d959dfe ;
    memory[2026] = 32'h3de776a5 ;
    memory[2027] = 32'hbe2091a6 ;
    memory[2028] = 32'hbbe72a8b ;
    memory[2029] = 32'hbdab6598 ;
    memory[2030] = 32'h3c966e75 ;
    memory[2031] = 32'hbcb8f94c ;
    memory[2032] = 32'hbdb665a9 ;
    memory[2033] = 32'hbd6f3bbe ;
    memory[2034] = 32'h3e0f2e75 ;
    memory[2035] = 32'h3d95dc87 ;
    memory[2036] = 32'hbe0bb8d3 ;
    memory[2037] = 32'hbe39845e ;
    memory[2038] = 32'h3d809301 ;
    memory[2039] = 32'h3dc79738 ;
    memory[2040] = 32'hbc34406d ;
    memory[2041] = 32'h3e064398 ;
    memory[2042] = 32'h3e120662 ;
    memory[2043] = 32'h3d0e6227 ;
    memory[2044] = 32'h3cd4a6ed ;
    memory[2045] = 32'hbe069392 ;
    memory[2046] = 32'h3e15279c ;
    memory[2047] = 32'hbdddfbc5 ;
    memory[2048] = 32'h3d7edaa3 ;
    memory[2049] = 32'h3e25b816 ;
    memory[2050] = 32'hbbc603ab ;
    memory[2051] = 32'h3d343d43 ;
    memory[2052] = 32'hbe1faff1 ;
    memory[2053] = 32'hbe1a95be ;
    memory[2054] = 32'hbbd69e5f ;
    memory[2055] = 32'hbbff4ec5 ;
    memory[2056] = 32'hbda6adab ;
    memory[2057] = 32'h3dba86ed ;
    memory[2058] = 32'hbdfd20ed ;
    memory[2059] = 32'h3dbab409 ;
    memory[2060] = 32'hbc94779f ;
    memory[2061] = 32'h3e30c300 ;
    memory[2062] = 32'h3d9212e0 ;
    memory[2063] = 32'h3d619037 ;
    memory[2064] = 32'h3dc4810a ;
    memory[2065] = 32'hbd3ffb6b ;
    memory[2066] = 32'hbbd0fb1c ;
    memory[2067] = 32'h3e23cb7f ;
    memory[2068] = 32'h3e2c846b ;
    memory[2069] = 32'h3ce2243e ;
    memory[2070] = 32'hbddac6d2 ;
    memory[2071] = 32'hbd0c612a ;
    memory[2072] = 32'h3d22b180 ;
    memory[2073] = 32'h3acd6e4b ;
    memory[2074] = 32'hbe2a4d26 ;
    memory[2075] = 32'h3e2f01c4 ;
    memory[2076] = 32'hbe111551 ;
    memory[2077] = 32'h3de24c57 ;
    memory[2078] = 32'hbd96a4de ;
    memory[2079] = 32'hbd82c5b6 ;
    memory[2080] = 32'h3e1d90c0 ;
    memory[2081] = 32'h3cd70289 ;
    memory[2082] = 32'h3d9236b3 ;
    memory[2083] = 32'h3c5deb76 ;
    memory[2084] = 32'h3c124896 ;
    memory[2085] = 32'hbd38fe4b ;
    memory[2086] = 32'h3c8fe895 ;
    memory[2087] = 32'h3c3bd685 ;
    memory[2088] = 32'hbdcb3535 ;
    memory[2089] = 32'h3cf80209 ;
    memory[2090] = 32'h3db0e212 ;
    memory[2091] = 32'h3e010477 ;
    memory[2092] = 32'h3b154f56 ;
    memory[2093] = 32'hbd9d19b1 ;
    memory[2094] = 32'hbdb86bc3 ;
    memory[2095] = 32'hbddbc0e0 ;
    memory[2096] = 32'hbe050f91 ;
    memory[2097] = 32'h3e2da14e ;
    memory[2098] = 32'hbdbc507e ;
    memory[2099] = 32'hbe19e8f1 ;
    memory[2100] = 32'hbdf3decc ;
    memory[2101] = 32'h3c541755 ;
    memory[2102] = 32'hbe3b8ff3 ;
    memory[2103] = 32'hbd27373e ;
    memory[2104] = 32'hbe1436d8 ;
    memory[2105] = 32'h3be82bf5 ;
    memory[2106] = 32'h3d77a169 ;
    memory[2107] = 32'h3d57c990 ;
    memory[2108] = 32'hbdff637c ;
    memory[2109] = 32'hbdc78d96 ;
    memory[2110] = 32'hbdfca78c ;
    memory[2111] = 32'h3d1cf6f2 ;
    memory[2112] = 32'hbe178012 ;
    memory[2113] = 32'h3e2d2c76 ;
    memory[2114] = 32'hbce6ded6 ;
    memory[2115] = 32'hba837416 ;
    memory[2116] = 32'h3dcd909e ;
    memory[2117] = 32'h3e3d41d0 ;
    memory[2118] = 32'h3de97cee ;
    memory[2119] = 32'h3dfea6ba ;
    memory[2120] = 32'h3de312f5 ;
    memory[2121] = 32'hbc5d9116 ;
    memory[2122] = 32'h3d81d105 ;
    memory[2123] = 32'h3df36775 ;
    memory[2124] = 32'h3e08b9b2 ;
    memory[2125] = 32'h3c90e8f0 ;
    memory[2126] = 32'hbd3c75d7 ;
    memory[2127] = 32'h3c34b9cd ;
    memory[2128] = 32'h3dc3f7c8 ;
    memory[2129] = 32'hbd65314c ;
    memory[2130] = 32'h3e0dba67 ;
    memory[2131] = 32'hbabe2018 ;
    memory[2132] = 32'hbe1c622f ;
    memory[2133] = 32'hbdd3da64 ;
    memory[2134] = 32'hbd99ff5f ;
    memory[2135] = 32'h3d682055 ;
    memory[2136] = 32'hbca13fc8 ;
    memory[2137] = 32'hbe0e854e ;
    memory[2138] = 32'hbdc04ed9 ;
    memory[2139] = 32'h3d40f158 ;
    memory[2140] = 32'hbc7fcb13 ;
    memory[2141] = 32'hbc8093f7 ;
    memory[2142] = 32'hbe1ba267 ;
    memory[2143] = 32'h3d32e6d8 ;
    memory[2144] = 32'h3e0ab67a ;
    memory[2145] = 32'hbd259650 ;
    memory[2146] = 32'hbd61b7eb ;
    memory[2147] = 32'hbe090cae ;
    memory[2148] = 32'h3c95d022 ;
    memory[2149] = 32'hbe177561 ;
    memory[2150] = 32'hbdb35d0a ;
    memory[2151] = 32'hbe172ffa ;
    memory[2152] = 32'hbe02b732 ;
    memory[2153] = 32'hbd091b80 ;
    memory[2154] = 32'hbd8f45b2 ;
    memory[2155] = 32'h3c61f33c ;
    memory[2156] = 32'hbd7c5ed6 ;
    memory[2157] = 32'hbc188ec7 ;
    memory[2158] = 32'hbd8cbaee ;
    memory[2159] = 32'h3cd28159 ;
    memory[2160] = 32'hbe4e9b9a ;
    memory[2161] = 32'hbda6f4cc ;
    memory[2162] = 32'hbe21c3e5 ;
    memory[2163] = 32'h3c862f26 ;
    memory[2164] = 32'h3cfdff03 ;
    memory[2165] = 32'h3d05dd48 ;
    memory[2166] = 32'hbcea7e0d ;
    memory[2167] = 32'h3d98fd4e ;
    memory[2168] = 32'hbe3a3dde ;
    memory[2169] = 32'hbddbd473 ;
    memory[2170] = 32'h3d0cb49a ;
    memory[2171] = 32'h3e012a12 ;
    memory[2172] = 32'h3df2e305 ;
    memory[2173] = 32'hbe48f8b6 ;
    memory[2174] = 32'h3e2bf0b8 ;
    memory[2175] = 32'hbd9c87cb ;
    memory[2176] = 32'h3e387777 ;
    memory[2177] = 32'hbd417eef ;
    memory[2178] = 32'h3e060b1c ;
    memory[2179] = 32'hbd951159 ;
    memory[2180] = 32'hbd8d7736 ;
    memory[2181] = 32'h3df96f44 ;
    memory[2182] = 32'hbdca62b6 ;
    memory[2183] = 32'hbd9cc651 ;
    memory[2184] = 32'hbe27b0c5 ;
    memory[2185] = 32'hbdd92544 ;
    memory[2186] = 32'h3daa44b2 ;
    memory[2187] = 32'h3e20f9e5 ;
    memory[2188] = 32'hbd7285ed ;
    memory[2189] = 32'h3dd50b27 ;
    memory[2190] = 32'h3dae024d ;
    memory[2191] = 32'hbcb94816 ;
    memory[2192] = 32'h3df8a4d2 ;
    memory[2193] = 32'hbdfffabb ;
    memory[2194] = 32'h3cbc44f1 ;
    memory[2195] = 32'hbde55ac4 ;
    memory[2196] = 32'h3d9126ea ;
    memory[2197] = 32'hbdb01125 ;
    memory[2198] = 32'h3d768854 ;
    memory[2199] = 32'hbe0534cd ;
    memory[2200] = 32'hbdba0f3b ;
    memory[2201] = 32'h3d394c43 ;
    memory[2202] = 32'hbc76ff47 ;
    memory[2203] = 32'hbb233e4b ;
    memory[2204] = 32'hbe27083f ;
    memory[2205] = 32'h3d96b5c6 ;
    memory[2206] = 32'hbe5f74c7 ;
    memory[2207] = 32'h3c618374 ;
    memory[2208] = 32'h3e20caba ;
    memory[2209] = 32'h3da50886 ;
    memory[2210] = 32'h3e0107f5 ;
    memory[2211] = 32'hbd28e2e7 ;
    memory[2212] = 32'h3c950500 ;
    memory[2213] = 32'hbbd3cc56 ;
    memory[2214] = 32'hbd09c5ee ;
    memory[2215] = 32'h3d11ed72 ;
    memory[2216] = 32'hbe0ad3da ;
    memory[2217] = 32'hbe20fc2c ;
    memory[2218] = 32'hbdeddb6a ;
    memory[2219] = 32'hbdfbe506 ;
    memory[2220] = 32'hbcacdab9 ;
    memory[2221] = 32'hbe0aeb0b ;
    memory[2222] = 32'h3ce546f3 ;
    memory[2223] = 32'hbbf989f7 ;
    memory[2224] = 32'h3dee1dd3 ;
    memory[2225] = 32'hbccc6197 ;
    memory[2226] = 32'hbddd0aa4 ;
    memory[2227] = 32'h3d2ad023 ;
    memory[2228] = 32'hbe3cff0e ;
    memory[2229] = 32'hbd02d073 ;
    memory[2230] = 32'hbe08067b ;
    memory[2231] = 32'h3e14e22c ;
    memory[2232] = 32'h3dc0da4f ;
    memory[2233] = 32'hbdb8dae3 ;
    memory[2234] = 32'hbe165918 ;
    memory[2235] = 32'hbd9396c2 ;
    memory[2236] = 32'h3c04dec8 ;
    memory[2237] = 32'hbdde636b ;
    memory[2238] = 32'h3d0df8d1 ;
    memory[2239] = 32'h3e06d653 ;
    memory[2240] = 32'hbba626b8 ;
    memory[2241] = 32'h3dc91dc3 ;
    memory[2242] = 32'hbe090454 ;
    memory[2243] = 32'hbd25e110 ;
    memory[2244] = 32'h3e1e3ab7 ;
    memory[2245] = 32'h3e2a934d ;
    memory[2246] = 32'h3d7c631e ;
    memory[2247] = 32'hbd2d9382 ;
    memory[2248] = 32'h3d0d9066 ;
    memory[2249] = 32'h3cf2260f ;
    memory[2250] = 32'hbe253df8 ;
    memory[2251] = 32'h3e15e279 ;
    memory[2252] = 32'hbdfe3d41 ;
    memory[2253] = 32'h3d79dc37 ;
    memory[2254] = 32'hbdd4cffa ;
    memory[2255] = 32'h3d8ee9b3 ;
    memory[2256] = 32'hbe003a5f ;
    memory[2257] = 32'h3e1abc0a ;
    memory[2258] = 32'hbd034b74 ;
    memory[2259] = 32'h3da82137 ;
    memory[2260] = 32'h3db0e757 ;
    memory[2261] = 32'h3e077950 ;
    memory[2262] = 32'h3d110058 ;
    memory[2263] = 32'h3da9cda0 ;
    memory[2264] = 32'hbbb2f0ce ;
    memory[2265] = 32'hbd62aadf ;
    memory[2266] = 32'h3ca836a0 ;
    memory[2267] = 32'hbc54e448 ;
    memory[2268] = 32'h39f526ac ;
    memory[2269] = 32'h3d751980 ;
    memory[2270] = 32'hbcb13c2d ;
    memory[2271] = 32'h3e2ef22c ;
    memory[2272] = 32'h3cb027c8 ;
    memory[2273] = 32'h3c7cd0c4 ;
    memory[2274] = 32'h3e15e6c6 ;
    memory[2275] = 32'h3e26216f ;
    memory[2276] = 32'hbdad4231 ;
    memory[2277] = 32'h3e05ccd5 ;
    memory[2278] = 32'h3a654c51 ;
    memory[2279] = 32'h3e2c707f ;
    memory[2280] = 32'h3e1c154e ;
    memory[2281] = 32'h3ced23fe ;
    memory[2282] = 32'hbd1c8f05 ;
    memory[2283] = 32'hbe1c774d ;
    memory[2284] = 32'hbde095eb ;
    memory[2285] = 32'h3db5c484 ;
    memory[2286] = 32'hbe21907a ;
    memory[2287] = 32'hbd916de3 ;
    memory[2288] = 32'h3ccef63d ;
    memory[2289] = 32'hbc10b3ff ;
    memory[2290] = 32'h3e06407c ;
    memory[2291] = 32'h3dc8249a ;
    memory[2292] = 32'hbe006979 ;
    memory[2293] = 32'hbd26c07a ;
    memory[2294] = 32'h3ccd20c8 ;
    memory[2295] = 32'h3df4921b ;
    memory[2296] = 32'hbd9adf91 ;
    memory[2297] = 32'h3e2e28b9 ;
    memory[2298] = 32'hbe0a4ec9 ;
    memory[2299] = 32'hbe05fa9c ;
    memory[2300] = 32'h3d417cc0 ;
    memory[2301] = 32'h3da93056 ;
    memory[2302] = 32'hbd18f867 ;
    memory[2303] = 32'h3e226590 ;
    memory[2304] = 32'h3e061a87 ;
    memory[2305] = 32'hbe2d86d4 ;
    memory[2306] = 32'h3e1239cb ;
    memory[2307] = 32'hbdc0d158 ;
    memory[2308] = 32'hbde26d82 ;
    memory[2309] = 32'h3e274a9d ;
    memory[2310] = 32'hbd602258 ;
    memory[2311] = 32'h3d74faa8 ;
    memory[2312] = 32'hbe29616a ;
    memory[2313] = 32'hbe1f3634 ;
    memory[2314] = 32'h3e52d9ea ;
    memory[2315] = 32'hbde2eee0 ;
    memory[2316] = 32'h3d306f41 ;
    memory[2317] = 32'h3e1f3c67 ;
    memory[2318] = 32'h3db5cf53 ;
    memory[2319] = 32'h3d5375ce ;
    memory[2320] = 32'hbd20ba0b ;
    memory[2321] = 32'h3c0968c8 ;
    memory[2322] = 32'hbdf5cc54 ;
    memory[2323] = 32'hbd833762 ;
    memory[2324] = 32'h3e02d576 ;
    memory[2325] = 32'hbd1b843c ;
    memory[2326] = 32'hbe3b9ec4 ;
    memory[2327] = 32'hbe169fb0 ;
    memory[2328] = 32'hbdeb9d53 ;
    memory[2329] = 32'hbd8f584d ;
    memory[2330] = 32'hbe219c15 ;
    memory[2331] = 32'hbe183a6c ;
    memory[2332] = 32'h3b9a36a7 ;
    memory[2333] = 32'h3c08959f ;
    memory[2334] = 32'h3e43bfd3 ;
    memory[2335] = 32'hbd01f221 ;
    memory[2336] = 32'h3dac3d25 ;
    memory[2337] = 32'hbe075a35 ;
    memory[2338] = 32'hbda68e9a ;
    memory[2339] = 32'h3db64b79 ;
    memory[2340] = 32'h3e100566 ;
    memory[2341] = 32'h3d135905 ;
    memory[2342] = 32'h3cebfce9 ;
    memory[2343] = 32'hbda14716 ;
    memory[2344] = 32'hbda6c45e ;
    memory[2345] = 32'hbbf67c26 ;
    memory[2346] = 32'hbc072857 ;
    memory[2347] = 32'h3d311f4d ;
    memory[2348] = 32'h3cc469c9 ;
    memory[2349] = 32'hbda6bf7d ;
    memory[2350] = 32'hbd8f4678 ;
    memory[2351] = 32'h3e3fca98 ;
    memory[2352] = 32'hbde6ac15 ;
    memory[2353] = 32'hbcdf6dbb ;
    memory[2354] = 32'hbdaecf9a ;
    memory[2355] = 32'hbde9a928 ;
    memory[2356] = 32'hbde1f854 ;
    memory[2357] = 32'hbe28e21d ;
    memory[2358] = 32'hbdf8726e ;
    memory[2359] = 32'h3d2217be ;
    memory[2360] = 32'h3d92c2e9 ;
    memory[2361] = 32'hbdaf95e2 ;
    memory[2362] = 32'h3e0f8742 ;
    memory[2363] = 32'hbdc898da ;
    memory[2364] = 32'h3e58b491 ;
    memory[2365] = 32'h3d89e96f ;
    memory[2366] = 32'hbd123258 ;
    memory[2367] = 32'h3d42a7db ;
    memory[2368] = 32'h3d8f2674 ;
    memory[2369] = 32'h3cf2bbdf ;
    memory[2370] = 32'hbe3dd028 ;
    memory[2371] = 32'hbe0995e4 ;
    memory[2372] = 32'hbe34118a ;
    memory[2373] = 32'hbe06d725 ;
    memory[2374] = 32'hbe2fc267 ;
    memory[2375] = 32'h3df23e0a ;
    memory[2376] = 32'hbe4e080f ;
    memory[2377] = 32'hbdf0bd1f ;
    memory[2378] = 32'h3e0833cc ;
    memory[2379] = 32'hbda75aad ;
    memory[2380] = 32'h3d0fb526 ;
    memory[2381] = 32'h3e16a9fd ;
    memory[2382] = 32'h3e29f08e ;
    memory[2383] = 32'h3da6676a ;
    memory[2384] = 32'hbe2d2685 ;
    memory[2385] = 32'h3dec6fc3 ;
    memory[2386] = 32'h3cdb11cf ;
    memory[2387] = 32'hbce4a920 ;
    memory[2388] = 32'hbd5fd869 ;
    memory[2389] = 32'hbcfe193f ;
    memory[2390] = 32'hbd17d685 ;
    memory[2391] = 32'hbd472a48 ;
    memory[2392] = 32'hbe39d785 ;
    memory[2393] = 32'hbb5944cf ;
    memory[2394] = 32'hbdd612f8 ;
    memory[2395] = 32'hbe372b9a ;
    memory[2396] = 32'h3d88416e ;
    memory[2397] = 32'h3df38a15 ;
    memory[2398] = 32'h3d0190ef ;
    memory[2399] = 32'hbdfa4d0a ;
    memory[2400] = 32'h3dc45cbb ;
    memory[2401] = 32'h3d1d105d ;
    memory[2402] = 32'hbe1b774f ;
    memory[2403] = 32'h3d2240a0 ;
    memory[2404] = 32'h3e2c08d5 ;
    memory[2405] = 32'h3dcd8d74 ;
    memory[2406] = 32'hbda5135f ;
    memory[2407] = 32'h3d77135f ;
    memory[2408] = 32'hbddb6491 ;
    memory[2409] = 32'hbe141988 ;
    memory[2410] = 32'hbd4a7783 ;
    memory[2411] = 32'h3bb67378 ;
    memory[2412] = 32'h3e242079 ;
    memory[2413] = 32'hbd8af1a0 ;
    memory[2414] = 32'h3e07d0fd ;
    memory[2415] = 32'hbd477d13 ;
    memory[2416] = 32'h3e2f8f75 ;
    memory[2417] = 32'hbde50fe0 ;
    memory[2418] = 32'h3e33b337 ;
    memory[2419] = 32'h3ce11a8f ;
    memory[2420] = 32'h3dbbfb1d ;
    memory[2421] = 32'hbd7d8755 ;
    memory[2422] = 32'h3d518547 ;
    memory[2423] = 32'h3c0e1ebc ;
    memory[2424] = 32'h3d00f3d7 ;
    memory[2425] = 32'hbe27de61 ;
    memory[2426] = 32'hbd0d5076 ;
    memory[2427] = 32'h3e39b396 ;
    memory[2428] = 32'h3e2a6a41 ;
    memory[2429] = 32'h3e04cdc1 ;
    memory[2430] = 32'hba946118 ;
    memory[2431] = 32'h3e013247 ;
    memory[2432] = 32'h3d78cc37 ;
    memory[2433] = 32'hbe18b272 ;
    memory[2434] = 32'hbdd4f76b ;
    memory[2435] = 32'h3d5300f5 ;
    memory[2436] = 32'hbd9200cf ;
    memory[2437] = 32'hbdfdc903 ;
    memory[2438] = 32'h3e1e458e ;
    memory[2439] = 32'hbe2e3e67 ;
    memory[2440] = 32'hbdc7fa14 ;
    memory[2441] = 32'h3dacefbd ;
    memory[2442] = 32'h3db9b837 ;
    memory[2443] = 32'h3e231947 ;
    memory[2444] = 32'h3d8775a9 ;
    memory[2445] = 32'hbdd0dca8 ;
    memory[2446] = 32'hbdf1ae3a ;
    memory[2447] = 32'hbe23d081 ;
    memory[2448] = 32'hbc9dec39 ;
    memory[2449] = 32'hbe0aac0e ;
    memory[2450] = 32'h3d9f341e ;
    memory[2451] = 32'hbe1e133d ;
    memory[2452] = 32'h3d11a6c2 ;
    memory[2453] = 32'hbde6f88e ;
    memory[2454] = 32'h3dbd3ee2 ;
    memory[2455] = 32'hbd866749 ;
    memory[2456] = 32'hbd3f21df ;
    memory[2457] = 32'hbc9f943d ;
    memory[2458] = 32'h3c9f57e8 ;
    memory[2459] = 32'h3d313e7c ;
    memory[2460] = 32'hbdf2c336 ;
    memory[2461] = 32'hbdb6c04c ;
    memory[2462] = 32'hbc5786e7 ;
    memory[2463] = 32'hbbe46d66 ;
    memory[2464] = 32'hbe037a1d ;
    memory[2465] = 32'hbe13f2a4 ;
    memory[2466] = 32'hbe21ff53 ;
    memory[2467] = 32'hbe03f414 ;
    memory[2468] = 32'h3e26cdfe ;
    memory[2469] = 32'hbd949586 ;
    memory[2470] = 32'hbbacf68b ;
    memory[2471] = 32'hbda4f1fa ;
    memory[2472] = 32'hbe2c0652 ;
    memory[2473] = 32'hbe0c3d2d ;
    memory[2474] = 32'h3dea3346 ;
    memory[2475] = 32'hbd20e7de ;
    memory[2476] = 32'hbb86822c ;
    memory[2477] = 32'h3a78de8c ;
    memory[2478] = 32'hbad225e6 ;
    memory[2479] = 32'hbdf3606d ;
    memory[2480] = 32'hbd089d08 ;
    memory[2481] = 32'hbe0f659e ;
    memory[2482] = 32'h3ddd5bf4 ;
    memory[2483] = 32'h3db9aacb ;
    memory[2484] = 32'h3e372147 ;
    memory[2485] = 32'hbde328b6 ;
    memory[2486] = 32'hbd35a566 ;
    memory[2487] = 32'h3d9a4d13 ;
    memory[2488] = 32'hbd192f7c ;
    memory[2489] = 32'h3d3052ed ;
    memory[2490] = 32'h3d9b8dc5 ;
    memory[2491] = 32'h3a5b80c9 ;
    memory[2492] = 32'hbccb1311 ;
    memory[2493] = 32'h3e322650 ;
    memory[2494] = 32'h3e38413d ;
    memory[2495] = 32'h3d83eeb6 ;
    memory[2496] = 32'hbe4776b0 ;
    memory[2497] = 32'h3dedf8b3 ;
    memory[2498] = 32'hbe2876b2 ;
    memory[2499] = 32'h3e24b63f ;
    memory[2500] = 32'h3da84c27 ;
    memory[2501] = 32'hbe0042be ;
    memory[2502] = 32'hbdd0309d ;
    memory[2503] = 32'hbd461f17 ;
    memory[2504] = 32'h3c2ab533 ;
    memory[2505] = 32'hbc049069 ;
    memory[2506] = 32'hbddf8350 ;
    memory[2507] = 32'h3de7c554 ;
    memory[2508] = 32'h3d235e15 ;
    memory[2509] = 32'h3d526103 ;
    memory[2510] = 32'hbe040ef7 ;
    memory[2511] = 32'h3e1802a4 ;
    memory[2512] = 32'h3e166d8e ;
    memory[2513] = 32'hbe06f6ec ;
    memory[2514] = 32'hbd9449c6 ;
    memory[2515] = 32'hbd2cedb8 ;
    memory[2516] = 32'h3d8ad205 ;
    memory[2517] = 32'h3df3c62f ;
    memory[2518] = 32'h3ca10799 ;
    memory[2519] = 32'hbdb9e25e ;
    memory[2520] = 32'h3e0f104f ;
    memory[2521] = 32'hbe6252f7 ;
    memory[2522] = 32'h3dea0e51 ;
    memory[2523] = 32'h3d1db2b4 ;
    memory[2524] = 32'h3dcd1294 ;
    memory[2525] = 32'h3d16ace6 ;
    memory[2526] = 32'h3d660c33 ;
    memory[2527] = 32'h3e1521f0 ;
    memory[2528] = 32'h3e1b2639 ;
    memory[2529] = 32'h3dcdf325 ;
    memory[2530] = 32'hbcaef570 ;
    memory[2531] = 32'hbb8525f6 ;
    memory[2532] = 32'hbd042b6b ;
    memory[2533] = 32'hbd637cb9 ;
    memory[2534] = 32'h3dd73d52 ;
    memory[2535] = 32'h3c62ad75 ;
    memory[2536] = 32'h3e19f637 ;
    memory[2537] = 32'h3e39f395 ;
    memory[2538] = 32'h3e2af760 ;
    memory[2539] = 32'h3e1ab824 ;
    memory[2540] = 32'hbcafdbde ;
    memory[2541] = 32'hbd64748f ;
    memory[2542] = 32'hbd4056fb ;
    memory[2543] = 32'hbe36aad7 ;
    memory[2544] = 32'h3ddb9065 ;
    memory[2545] = 32'h3dbc1c50 ;
    memory[2546] = 32'h3d3f7b42 ;
    memory[2547] = 32'h3d8703e6 ;
    memory[2548] = 32'h3c4ff6b2 ;
    memory[2549] = 32'h3d2afa18 ;
    memory[2550] = 32'hbe180d41 ;
    memory[2551] = 32'h3cf06b87 ;
    memory[2552] = 32'hbd921363 ;
    memory[2553] = 32'h3ce01de1 ;
    memory[2554] = 32'hbe1a6efc ;
    memory[2555] = 32'hbdcd0b44 ;
    memory[2556] = 32'h3cc052bd ;
    memory[2557] = 32'hbd55b582 ;
    memory[2558] = 32'hbd9ffa5c ;
    memory[2559] = 32'h3dc25c26 ;
    memory[2560] = 32'hbdabc38b ;
    memory[2561] = 32'hbb4fc6f8 ;
    memory[2562] = 32'hbde0324a ;
    memory[2563] = 32'hbd279fe2 ;
    memory[2564] = 32'h3d8a9f58 ;
    memory[2565] = 32'h3d4062ca ;
    memory[2566] = 32'h3d425a28 ;
    memory[2567] = 32'h3d6f3d6b ;
    memory[2568] = 32'hbd6b2a9f ;
    memory[2569] = 32'h3df5935e ;
    memory[2570] = 32'hbdefcb73 ;
    memory[2571] = 32'h3e2184d5 ;
    memory[2572] = 32'hbd8cb127 ;
    memory[2573] = 32'h3e18f0b0 ;
    memory[2574] = 32'h3dc72bf3 ;
    memory[2575] = 32'hbe18afd7 ;
    memory[2576] = 32'hbd7449bc ;
    memory[2577] = 32'hbd6eb6b4 ;
    memory[2578] = 32'hbe21d919 ;
    memory[2579] = 32'h3cc6eab2 ;
    memory[2580] = 32'hbda90b37 ;
    memory[2581] = 32'hbd0f8b72 ;
    memory[2582] = 32'hbd1987b2 ;
    memory[2583] = 32'hbd107f3a ;
    memory[2584] = 32'hbc9fe4b4 ;
    memory[2585] = 32'h3d845411 ;
    memory[2586] = 32'hbe003c54 ;
    memory[2587] = 32'h3d9f93e0 ;
    memory[2588] = 32'h3d21cf95 ;
    memory[2589] = 32'h3df1a378 ;
    memory[2590] = 32'hbe1bb588 ;
    memory[2591] = 32'h3e559819 ;
    memory[2592] = 32'h3df03599 ;
    memory[2593] = 32'hbda562a9 ;
    memory[2594] = 32'hbd69a926 ;
    memory[2595] = 32'h3e259ff8 ;
    memory[2596] = 32'h3bbd8f26 ;
    memory[2597] = 32'h3db41a20 ;
    memory[2598] = 32'hbc85bd75 ;
    memory[2599] = 32'h3d8cf860 ;
    memory[2600] = 32'hbce42d5a ;
    memory[2601] = 32'hbcfeef68 ;
    memory[2602] = 32'h3e0ac0bc ;
    memory[2603] = 32'hbdd83943 ;
    memory[2604] = 32'hbe23236f ;
    memory[2605] = 32'h3d48cff5 ;
    memory[2606] = 32'hbdcad149 ;
    memory[2607] = 32'h3d9bbea7 ;
    memory[2608] = 32'hbdb9cefc ;
    memory[2609] = 32'hbe0f0b7b ;
    memory[2610] = 32'h3e0fd6fd ;
    memory[2611] = 32'h3d1a285e ;
    memory[2612] = 32'hbd446934 ;
    memory[2613] = 32'hbdd27b2b ;
    memory[2614] = 32'hbd890468 ;
    memory[2615] = 32'hbe015d77 ;
    memory[2616] = 32'hbe0b5a1e ;
    memory[2617] = 32'h3d447c79 ;
    memory[2618] = 32'hbd57a749 ;
    memory[2619] = 32'hbd8559ea ;
    memory[2620] = 32'h3cb463de ;
    memory[2621] = 32'hbe28bc30 ;
    memory[2622] = 32'h3d0021e4 ;
    memory[2623] = 32'hbcfb9ec6 ;
    memory[2624] = 32'hbdc62e8a ;
    memory[2625] = 32'h3d90fa69 ;
    memory[2626] = 32'hbe5999bc ;
    memory[2627] = 32'h3cf01eb5 ;
    memory[2628] = 32'hbe0a1d27 ;
    memory[2629] = 32'h3da7df3d ;
    memory[2630] = 32'h3e1570ec ;
    memory[2631] = 32'hbda839ae ;
    memory[2632] = 32'h389b0201 ;
    memory[2633] = 32'hbdc91d39 ;
    memory[2634] = 32'hbe16f2bd ;
    memory[2635] = 32'h3d835551 ;
    memory[2636] = 32'hbdc658dd ;
    memory[2637] = 32'hbe391918 ;
    memory[2638] = 32'h3defd178 ;
    memory[2639] = 32'hbc8cff9c ;
    memory[2640] = 32'h3dc85237 ;
    memory[2641] = 32'h3e089620 ;
    memory[2642] = 32'h3db79cd8 ;
    memory[2643] = 32'hbd9ab6cd ;
    memory[2644] = 32'hbd27dabc ;
    memory[2645] = 32'h3d133996 ;
    memory[2646] = 32'h3e363a8c ;
    memory[2647] = 32'h3dee206a ;
    memory[2648] = 32'h3d7d0cd7 ;
    memory[2649] = 32'h3e3bd7b0 ;
    memory[2650] = 32'h3e2f4053 ;
    memory[2651] = 32'hbcc3ec32 ;
    memory[2652] = 32'hbe004a53 ;
    memory[2653] = 32'hbcf5abcc ;
    memory[2654] = 32'h3d239112 ;
    memory[2655] = 32'h3e40d28c ;
    memory[2656] = 32'hbd0e5ab7 ;
    memory[2657] = 32'h3d330de7 ;
    memory[2658] = 32'h3d549a61 ;
    memory[2659] = 32'h3e223a8e ;
    memory[2660] = 32'h3c9f823e ;
    memory[2661] = 32'hbd6b9b1b ;
    memory[2662] = 32'hbde3e8f6 ;
    memory[2663] = 32'hbd9e07e3 ;
    memory[2664] = 32'hbe1f4e30 ;
    memory[2665] = 32'hbe366895 ;
    memory[2666] = 32'h3daa511a ;
    memory[2667] = 32'hbdf4913a ;
    memory[2668] = 32'hbe006c58 ;
    memory[2669] = 32'hbd9be707 ;
    memory[2670] = 32'hbd272eb8 ;
    memory[2671] = 32'h3dc7ebf1 ;
    memory[2672] = 32'h3da06437 ;
    memory[2673] = 32'h3e481a9a ;
    memory[2674] = 32'hbe1a986a ;
    memory[2675] = 32'hbd1ee375 ;
    memory[2676] = 32'h3dd7efb0 ;
    memory[2677] = 32'h3e123349 ;
    memory[2678] = 32'h3da5fb73 ;
    memory[2679] = 32'h3e29af95 ;
    memory[2680] = 32'h3e2dfc98 ;
    memory[2681] = 32'hbd4af608 ;
    memory[2682] = 32'h3d55c3e0 ;
    memory[2683] = 32'h3e01d576 ;
    memory[2684] = 32'h3e167f9e ;
    memory[2685] = 32'h3e03b734 ;
    memory[2686] = 32'hbe3561d8 ;
    memory[2687] = 32'hbc3489a8 ;
    memory[2688] = 32'h3e299713 ;
    memory[2689] = 32'hbde8d277 ;
    memory[2690] = 32'h3d144643 ;
    memory[2691] = 32'hbd1dab4a ;
    memory[2692] = 32'h3dcecf0a ;
    memory[2693] = 32'hbd7c74a4 ;
    memory[2694] = 32'hbe1606e3 ;
    memory[2695] = 32'hbe15ef5b ;
    memory[2696] = 32'h3cfc7767 ;
    memory[2697] = 32'h3dde5809 ;
    memory[2698] = 32'hbd42db1f ;
    memory[2699] = 32'h3d750bf3 ;
    memory[2700] = 32'hbdf5f650 ;
    memory[2701] = 32'hbd159578 ;
    memory[2702] = 32'h3dd46cdc ;
    memory[2703] = 32'h3e3695ea ;
    memory[2704] = 32'h3dacdd25 ;
    memory[2705] = 32'h3b1c6ad9 ;
    memory[2706] = 32'h3e0d6189 ;
    memory[2707] = 32'h3da02568 ;
    memory[2708] = 32'hbdaf0c99 ;
    memory[2709] = 32'hbe06912d ;
    memory[2710] = 32'h3e22f60f ;
    memory[2711] = 32'h3ccf7774 ;
    memory[2712] = 32'hbc0e0d2a ;
    memory[2713] = 32'h3e2bc65b ;
    memory[2714] = 32'hbd7ed3a7 ;
    memory[2715] = 32'h3d5b2050 ;
    memory[2716] = 32'hbd8953c2 ;
    memory[2717] = 32'h3d70bad7 ;
    memory[2718] = 32'hbe13c2b5 ;
    memory[2719] = 32'hbda37906 ;
    memory[2720] = 32'hbdfe540b ;
    memory[2721] = 32'hbdd48749 ;
    memory[2722] = 32'hbd0db9da ;
    memory[2723] = 32'hbe2d567d ;
    memory[2724] = 32'h3dbcb0fb ;
    memory[2725] = 32'h3cebfc12 ;
    memory[2726] = 32'hbcd874dd ;
    memory[2727] = 32'h3d5729df ;
    memory[2728] = 32'hbe16b641 ;
    memory[2729] = 32'hbe055036 ;
    memory[2730] = 32'hbd9a1bf3 ;
    memory[2731] = 32'h3e0dc813 ;
    memory[2732] = 32'hbd564d40 ;
    memory[2733] = 32'h3cb35825 ;
    memory[2734] = 32'h3ddc143f ;
    memory[2735] = 32'h3dcb0a67 ;
    memory[2736] = 32'h3decd186 ;
    memory[2737] = 32'h3c9fb9c1 ;
    memory[2738] = 32'hbd7072e0 ;
    memory[2739] = 32'hbd663ea1 ;
    memory[2740] = 32'hbe1cac42 ;
    memory[2741] = 32'h3c452a98 ;
    memory[2742] = 32'hbd3438da ;
    memory[2743] = 32'hbb4feef9 ;
    memory[2744] = 32'h3d996125 ;
    memory[2745] = 32'h3e1ae8c6 ;
    memory[2746] = 32'hbe1a088b ;
    memory[2747] = 32'h3de68968 ;
    memory[2748] = 32'h3dd71ff4 ;
    memory[2749] = 32'hbcbefc30 ;
    memory[2750] = 32'h3d2fef79 ;
    memory[2751] = 32'hbe00d800 ;
    memory[2752] = 32'h3dd78221 ;
    memory[2753] = 32'h3d974028 ;
    memory[2754] = 32'hbd390749 ;
    memory[2755] = 32'h3d3b5c3f ;
    memory[2756] = 32'hbd6d21a8 ;
    memory[2757] = 32'hbd8e0783 ;
    memory[2758] = 32'hbdababaf ;
    memory[2759] = 32'hbde0c4ee ;
    memory[2760] = 32'hbdbb86c1 ;
    memory[2761] = 32'hbd1b2c0d ;
    memory[2762] = 32'hbd6521b7 ;
    memory[2763] = 32'hbd654bb5 ;
    memory[2764] = 32'h3e3441cf ;
    memory[2765] = 32'hbe37bbb2 ;
    memory[2766] = 32'h3d9232e1 ;
    memory[2767] = 32'h3e20629e ;
    memory[2768] = 32'h3e07a8f1 ;
    memory[2769] = 32'h3dd60664 ;
    memory[2770] = 32'h3dc811f6 ;
    memory[2771] = 32'h3daa3147 ;
    memory[2772] = 32'hbcce1e8f ;
    memory[2773] = 32'hbe1e9cc0 ;
    memory[2774] = 32'h3d158a05 ;
    memory[2775] = 32'hbe1e0dd8 ;
    memory[2776] = 32'h3c99633c ;
    memory[2777] = 32'h3dd00e2f ;
    memory[2778] = 32'h3d85989c ;
    memory[2779] = 32'h3e1ae844 ;
    memory[2780] = 32'h3db9f51b ;
    memory[2781] = 32'h3dab0741 ;
    memory[2782] = 32'hbe099d4d ;
    memory[2783] = 32'hbdb7f2a8 ;
    memory[2784] = 32'h3de57d57 ;
    memory[2785] = 32'h3e15038d ;
    memory[2786] = 32'hbe39b725 ;
    memory[2787] = 32'hbb523538 ;
    memory[2788] = 32'h3d56aea9 ;
    memory[2789] = 32'h3caead55 ;
    memory[2790] = 32'h3da1006f ;
    memory[2791] = 32'h3c33abc6 ;
    memory[2792] = 32'hbe354c42 ;
    memory[2793] = 32'hbe068aeb ;
    memory[2794] = 32'hbe086ca0 ;
    memory[2795] = 32'hbe197c95 ;
    memory[2796] = 32'h3dd49742 ;
    memory[2797] = 32'h3ceea035 ;
    memory[2798] = 32'h3c23b932 ;
    memory[2799] = 32'hbd0c9d8f ;
    memory[2800] = 32'hbce73dfe ;
    memory[2801] = 32'h3d09a573 ;
    memory[2802] = 32'hbd999c4f ;
    memory[2803] = 32'hbe123255 ;
    memory[2804] = 32'hbae466b7 ;
    memory[2805] = 32'h3ca4161a ;
    memory[2806] = 32'h3a9eb484 ;
    memory[2807] = 32'hbc6157a6 ;
    memory[2808] = 32'hbe08781e ;
    memory[2809] = 32'h3c12ba85 ;
    memory[2810] = 32'h3dd83a49 ;
    memory[2811] = 32'hbe2bf73d ;
    memory[2812] = 32'h3d8cac28 ;
    memory[2813] = 32'h3d6ddcb3 ;
    memory[2814] = 32'hbe254f2d ;
    memory[2815] = 32'hbe1cfb7b ;
    memory[2816] = 32'hbe36f7f4 ;
    memory[2817] = 32'h3db46be4 ;
    memory[2818] = 32'h3e0e686b ;
    memory[2819] = 32'hbdd8bb15 ;
    memory[2820] = 32'h3dc9759b ;
    memory[2821] = 32'hbe2ea35d ;
    memory[2822] = 32'hbd959b4a ;
    memory[2823] = 32'hbe31fc3f ;
    memory[2824] = 32'h3e0451b6 ;
    memory[2825] = 32'h3ddf2ed6 ;
    memory[2826] = 32'hbc93b9e9 ;
    memory[2827] = 32'h3e1f4443 ;
    memory[2828] = 32'h3de89fb9 ;
    memory[2829] = 32'h3c0b40a1 ;
    memory[2830] = 32'h3da8701b ;
    memory[2831] = 32'hbdeda792 ;
    memory[2832] = 32'h3e020a0a ;
    memory[2833] = 32'h3e1bd557 ;
    memory[2834] = 32'hbcbc698c ;
    memory[2835] = 32'h3db15e5a ;
    memory[2836] = 32'h3da89ebd ;
    memory[2837] = 32'hbccc7dd5 ;
    memory[2838] = 32'h3e4607b1 ;
    memory[2839] = 32'h3a53ebf9 ;
    memory[2840] = 32'h3cdae877 ;
    memory[2841] = 32'h3d0b2f24 ;
    memory[2842] = 32'h3db3a153 ;
    memory[2843] = 32'h3d94ef0b ;
    memory[2844] = 32'h3deb906a ;
    memory[2845] = 32'hbd42fccc ;
    memory[2846] = 32'h3ad9752f ;
    memory[2847] = 32'hbdae2dde ;
    memory[2848] = 32'hbd418775 ;
    memory[2849] = 32'hbdd01cb4 ;
    memory[2850] = 32'h3dbf3b75 ;
    memory[2851] = 32'h3e4ba091 ;
    memory[2852] = 32'hbd8f8391 ;
    memory[2853] = 32'hbe23f4db ;
    memory[2854] = 32'hbe075593 ;
    memory[2855] = 32'hbdfd54fa ;
    memory[2856] = 32'hbde147ed ;
    memory[2857] = 32'hbe0a8178 ;
    memory[2858] = 32'h3cbeb40b ;
    memory[2859] = 32'h3d5aa86e ;
    memory[2860] = 32'hbdbacd37 ;
    memory[2861] = 32'hbc50c3b5 ;
    memory[2862] = 32'h3e2d2c8a ;
    memory[2863] = 32'hbdb8ba5c ;
    memory[2864] = 32'h3dff99b1 ;
    memory[2865] = 32'h3e0d94bf ;
    memory[2866] = 32'h3e024b04 ;
    memory[2867] = 32'hbb0c0c9a ;
    memory[2868] = 32'hbd9d7784 ;
    memory[2869] = 32'hbd750ff9 ;
    memory[2870] = 32'hbd952580 ;
    memory[2871] = 32'h3e21c7a5 ;
    memory[2872] = 32'h3dfe3aa9 ;
    memory[2873] = 32'hbd9854b4 ;
    memory[2874] = 32'hbd683f44 ;
    memory[2875] = 32'hbd836b9b ;
    memory[2876] = 32'h3cf085f9 ;
    memory[2877] = 32'h3da453a9 ;
    memory[2878] = 32'h3c7e524e ;
    memory[2879] = 32'h3d2fbb0d ;
    memory[2880] = 32'h3cf7ea43 ;
    memory[2881] = 32'hbe1bc86a ;
    memory[2882] = 32'h3e1aefe9 ;
    memory[2883] = 32'h3e28ff20 ;
    memory[2884] = 32'h3cda0aea ;
    memory[2885] = 32'h3e37f753 ;
    memory[2886] = 32'hbdfc815a ;
    memory[2887] = 32'hbbbf61cd ;
    memory[2888] = 32'hbbee5408 ;
    memory[2889] = 32'h3e07535b ;
    memory[2890] = 32'hbd4b781e ;
    memory[2891] = 32'hbe28543b ;
    memory[2892] = 32'hbc2f7772 ;
    memory[2893] = 32'h3e182a1b ;
    memory[2894] = 32'h3e3445b4 ;
    memory[2895] = 32'hbd599af5 ;
    memory[2896] = 32'hbc29f8ad ;
    memory[2897] = 32'h3e1fc9fb ;
    memory[2898] = 32'hbe2a376b ;
    memory[2899] = 32'hbd781bc0 ;
    memory[2900] = 32'h3c6982f8 ;
    memory[2901] = 32'h3d9bd0de ;
    memory[2902] = 32'hbd83237f ;
    memory[2903] = 32'h3d94ad1f ;
    memory[2904] = 32'hbdae3535 ;
    memory[2905] = 32'h3d9f205e ;
    memory[2906] = 32'h3dfa0d44 ;
    memory[2907] = 32'hbe47ab91 ;
    memory[2908] = 32'hbe117e97 ;
    memory[2909] = 32'hbc911576 ;
    memory[2910] = 32'hbc98bbd2 ;
    memory[2911] = 32'h3e0b70c6 ;
    memory[2912] = 32'h3ca0c3a2 ;
    memory[2913] = 32'hbc54d32a ;
    memory[2914] = 32'hbbe7d5b8 ;
    memory[2915] = 32'hbdf8a65d ;
    memory[2916] = 32'hbe159583 ;
    memory[2917] = 32'h3ce3413d ;
    memory[2918] = 32'h3dd49c64 ;
    memory[2919] = 32'h3c0128a2 ;
    memory[2920] = 32'h3c77e4e9 ;
    memory[2921] = 32'h3c58f6dd ;
    memory[2922] = 32'h3e4ca4d0 ;
    memory[2923] = 32'hbd1cf81e ;
    memory[2924] = 32'hbd835f5c ;
    memory[2925] = 32'h3daec489 ;
    memory[2926] = 32'h3dc22710 ;
    memory[2927] = 32'hbd6c7299 ;
    memory[2928] = 32'hbe1ad1dd ;
    memory[2929] = 32'hbdb8e8c7 ;
    memory[2930] = 32'h3d1933d1 ;
    memory[2931] = 32'h3c91b948 ;
    memory[2932] = 32'h3e462277 ;
    memory[2933] = 32'hbdc09d6a ;
    memory[2934] = 32'h3d9939f5 ;
    memory[2935] = 32'h3de03f94 ;
    memory[2936] = 32'h3ddd5dc8 ;
    memory[2937] = 32'hbe3fb086 ;
    memory[2938] = 32'hbda74ea9 ;
    memory[2939] = 32'hbd8628f6 ;
    memory[2940] = 32'h3d69634c ;
    memory[2941] = 32'h3bba1f3c ;
    memory[2942] = 32'hbdfb95f2 ;
    memory[2943] = 32'hbc5399b5 ;
    memory[2944] = 32'hbd121a15 ;
    memory[2945] = 32'h3c2bf941 ;
    memory[2946] = 32'hbe2f99b3 ;
    memory[2947] = 32'hbc8deb1d ;
    memory[2948] = 32'h3e30a952 ;
    memory[2949] = 32'hbd877e86 ;
    memory[2950] = 32'h3d14986c ;
    memory[2951] = 32'hbe11c06d ;
    memory[2952] = 32'hbe4637e7 ;
    memory[2953] = 32'h3d3ec06a ;
    memory[2954] = 32'h3e028f9e ;
    memory[2955] = 32'hbe0eb506 ;
    memory[2956] = 32'hbda48ffa ;
    memory[2957] = 32'hbe02cf9e ;
    memory[2958] = 32'hbd67043e ;
    memory[2959] = 32'hbd879286 ;
    memory[2960] = 32'h3dc5128a ;
    memory[2961] = 32'hbd975f72 ;
    memory[2962] = 32'h3ca7813c ;
    memory[2963] = 32'hbd382298 ;
    memory[2964] = 32'h3e09ecb8 ;
    memory[2965] = 32'hbd00ec2f ;
    memory[2966] = 32'hbd82b7a0 ;
    memory[2967] = 32'h3e0c0937 ;
    memory[2968] = 32'hbd5e96cb ;
    memory[2969] = 32'hbe43e0f0 ;
    memory[2970] = 32'h3deac300 ;
    memory[2971] = 32'h3e36995e ;
    memory[2972] = 32'h3e08f470 ;
    memory[2973] = 32'hbd97afc3 ;
    memory[2974] = 32'h3ca08c8a ;
    memory[2975] = 32'hbdc8d139 ;
    memory[2976] = 32'h3d83bded ;
    memory[2977] = 32'h3e282ba3 ;
    memory[2978] = 32'h3d05633d ;
    memory[2979] = 32'h3dba6593 ;
    memory[2980] = 32'h3d89f296 ;
    memory[2981] = 32'h3c92c409 ;
    memory[2982] = 32'h3e1f03e1 ;
    memory[2983] = 32'hbcadbb67 ;
    memory[2984] = 32'h3db373f5 ;
    memory[2985] = 32'h3dcb7b2a ;
    memory[2986] = 32'hbdf13747 ;
    memory[2987] = 32'hbdfe963f ;
    memory[2988] = 32'hbd2b6b10 ;
    memory[2989] = 32'hbd3c1b8f ;
    memory[2990] = 32'h3c9a8ef9 ;
    memory[2991] = 32'h3d8810c9 ;
    memory[2992] = 32'h3ce3b13d ;
    memory[2993] = 32'hbe055fd0 ;
    memory[2994] = 32'h3db26ff3 ;
    memory[2995] = 32'h3d0b21a1 ;
    memory[2996] = 32'hbdcc4efb ;
    memory[2997] = 32'hbe22da30 ;
    memory[2998] = 32'hbc035b84 ;
    memory[2999] = 32'h3ca14c6b ;
    memory[3000] = 32'hbe0bf727 ;
    memory[3001] = 32'hbd016c9c ;
    memory[3002] = 32'hbd13efed ;
    memory[3003] = 32'hbdcfcfb9 ;
    memory[3004] = 32'hbdcf09ac ;
    memory[3005] = 32'hbdbf3ac7 ;
    memory[3006] = 32'hbd0559dc ;
    memory[3007] = 32'hbe20e0ce ;
    memory[3008] = 32'hbd836452 ;
    memory[3009] = 32'hbc1a4673 ;
    memory[3010] = 32'h3e2765b0 ;
    memory[3011] = 32'hbe283aa9 ;
    memory[3012] = 32'h3cca5e32 ;
    memory[3013] = 32'hbdc33b21 ;
    memory[3014] = 32'hba06b209 ;
    memory[3015] = 32'h3b97107b ;
    memory[3016] = 32'hbd21c176 ;
    memory[3017] = 32'h3dc07d8a ;
    memory[3018] = 32'hbdc76b5e ;
    memory[3019] = 32'hbdb60893 ;
    memory[3020] = 32'h3d623da2 ;
    memory[3021] = 32'h3d2c63e2 ;
    memory[3022] = 32'h3daeb080 ;
    memory[3023] = 32'h3db19b4c ;
    memory[3024] = 32'hbd82558e ;
    memory[3025] = 32'hbddc4dcd ;
    memory[3026] = 32'h3e13c8de ;
    memory[3027] = 32'h3dd6799b ;
    memory[3028] = 32'hbe42b818 ;
    memory[3029] = 32'hbe258f1d ;
    memory[3030] = 32'h3d1d1580 ;
    memory[3031] = 32'h3cc5906c ;
    memory[3032] = 32'hbdb059e9 ;
    memory[3033] = 32'hbce8e99a ;
    memory[3034] = 32'h3d6bfcc3 ;
    memory[3035] = 32'hbd653677 ;
    memory[3036] = 32'hbc97cec3 ;
    memory[3037] = 32'h3d409973 ;
    memory[3038] = 32'h3d641977 ;
    memory[3039] = 32'hbe067944 ;
    memory[3040] = 32'h3dac9b93 ;
    memory[3041] = 32'h3dce696b ;
    memory[3042] = 32'h3dc4a2ac ;
    memory[3043] = 32'h3b7ab1be ;
    memory[3044] = 32'h3dc7662f ;
    memory[3045] = 32'h3dc2e5e8 ;
    memory[3046] = 32'h3e16bbf7 ;
    memory[3047] = 32'hbd284877 ;
    memory[3048] = 32'h3e1c373f ;
    memory[3049] = 32'hbe3ae662 ;
    memory[3050] = 32'h3e1b70cf ;
    memory[3051] = 32'h3c6c6cb2 ;
    memory[3052] = 32'hbdc44b02 ;
    memory[3053] = 32'h3d47a8c4 ;
    memory[3054] = 32'hbd9b45a2 ;
    memory[3055] = 32'h3e1ce645 ;
    memory[3056] = 32'h3ba3c79e ;
    memory[3057] = 32'h3e3fae05 ;
    memory[3058] = 32'hbdcb3496 ;
    memory[3059] = 32'hbe365d10 ;
    memory[3060] = 32'hbe35e935 ;
    memory[3061] = 32'hbe01ac67 ;
    memory[3062] = 32'h3e0e547b ;
    memory[3063] = 32'hbd69ea18 ;
    memory[3064] = 32'hbd823ec1 ;
    memory[3065] = 32'h3c2bd54a ;
    memory[3066] = 32'h3d786384 ;
    memory[3067] = 32'hbd7bc4af ;
    memory[3068] = 32'hbe0c4a92 ;
    memory[3069] = 32'hbe44b9c7 ;
    memory[3070] = 32'h3d84df95 ;
    memory[3071] = 32'hbdcfee9d ;
    memory[3072] = 32'h3e046e3d ;
    memory[3073] = 32'h3d36be31 ;
    memory[3074] = 32'h3d923d16 ;
    memory[3075] = 32'h3df90937 ;
    memory[3076] = 32'hbdbc099c ;
    memory[3077] = 32'h3d9cf974 ;
    memory[3078] = 32'h3db65223 ;
    memory[3079] = 32'hba0f44b1 ;
    memory[3080] = 32'h3df3590c ;
    memory[3081] = 32'hbd5baaef ;
    memory[3082] = 32'h3cf0d753 ;
    memory[3083] = 32'hbda30a30 ;
    memory[3084] = 32'h3d2f4f52 ;
    memory[3085] = 32'hbe1cd855 ;
    memory[3086] = 32'hbe221313 ;
    memory[3087] = 32'h3d2a973f ;
    memory[3088] = 32'hbe1cc28b ;
    memory[3089] = 32'hbdd13115 ;
    memory[3090] = 32'h3dc4d3eb ;
    memory[3091] = 32'hbd4c8486 ;
    memory[3092] = 32'hbd480533 ;
    memory[3093] = 32'hbd566a4a ;
    memory[3094] = 32'hbdc7397e ;
    memory[3095] = 32'h3da12cad ;
    memory[3096] = 32'h3c7465be ;
    memory[3097] = 32'hbd1c972c ;
    memory[3098] = 32'hbe00fede ;
    memory[3099] = 32'hbd61992e ;
    memory[3100] = 32'h3d797cae ;
    memory[3101] = 32'h3e0b3d8b ;
    memory[3102] = 32'hbd0c8ebd ;
    memory[3103] = 32'hbda149a2 ;
    memory[3104] = 32'hbd7f7404 ;
    memory[3105] = 32'hbb6ebd71 ;
    memory[3106] = 32'h3d2875d2 ;
    memory[3107] = 32'hbe0372ae ;
    memory[3108] = 32'h3d606cb9 ;
    memory[3109] = 32'h3cd45665 ;
    memory[3110] = 32'h3d688ab8 ;
    memory[3111] = 32'hbdec2632 ;
    memory[3112] = 32'hbcb6e5d9 ;
    memory[3113] = 32'h3dd35e8d ;
    memory[3114] = 32'h3d47be02 ;
    memory[3115] = 32'hbd2d6006 ;
    memory[3116] = 32'hbd97eacc ;
    memory[3117] = 32'hbc9fc2a2 ;
    memory[3118] = 32'hbe118b51 ;
    memory[3119] = 32'hbdf13c22 ;
    memory[3120] = 32'hbe1af32b ;
    memory[3121] = 32'hbe0f7ec0 ;
    memory[3122] = 32'h3df74812 ;
    memory[3123] = 32'hbb6d7e7d ;
    memory[3124] = 32'h3d6a715e ;
    memory[3125] = 32'hbe05bab7 ;
    memory[3126] = 32'hbd22e863 ;
    memory[3127] = 32'h3d129c87 ;
    memory[3128] = 32'h3c20aaf6 ;
    memory[3129] = 32'hbe420ab7 ;
    memory[3130] = 32'h3ddab25c ;
    memory[3131] = 32'hbe17f731 ;
    memory[3132] = 32'hbd82ae88 ;
    memory[3133] = 32'h3dc5e601 ;
    memory[3134] = 32'hbd955d91 ;
    memory[3135] = 32'hbe049fe3 ;
    memory[3136] = 32'hbd3410a6 ;
    memory[3137] = 32'hbdaef57f ;
    memory[3138] = 32'h3c59c557 ;
    memory[3139] = 32'h3e22678f ;
    memory[3140] = 32'h3e12ec2e ;
    memory[3141] = 32'hbe2300a4 ;
    memory[3142] = 32'h3dedff0e ;
    memory[3143] = 32'h3e3f2198 ;
    memory[3144] = 32'hbd44a5e6 ;
    memory[3145] = 32'h3d9d59b7 ;
    memory[3146] = 32'h3e136e8e ;
    memory[3147] = 32'hbe0cf992 ;
    memory[3148] = 32'hbe189d32 ;
    memory[3149] = 32'hbd4d54bf ;
    memory[3150] = 32'hbe0dd2d9 ;
    memory[3151] = 32'h3dc41e13 ;
    memory[3152] = 32'h3d32425c ;
    memory[3153] = 32'hbccf29f9 ;
    memory[3154] = 32'hbdccc9d3 ;
    memory[3155] = 32'hbb21f79f ;
    memory[3156] = 32'h3e023f99 ;
    memory[3157] = 32'h3df9b9b5 ;
    memory[3158] = 32'h3e32bc79 ;
    memory[3159] = 32'hbe38c321 ;
    memory[3160] = 32'h3dd6060a ;
    memory[3161] = 32'h3c338451 ;
    memory[3162] = 32'hbe233c36 ;
    memory[3163] = 32'h3e16de4a ;
    memory[3164] = 32'h3de8a9da ;
    memory[3165] = 32'h3dfefad1 ;
    memory[3166] = 32'hbbf669d9 ;
    memory[3167] = 32'hbdd59b01 ;
    memory[3168] = 32'h3e1b5f28 ;
    memory[3169] = 32'hbe290832 ;
    memory[3170] = 32'h3c03d5dd ;
    memory[3171] = 32'hbde3f0de ;
    memory[3172] = 32'hbdbc3913 ;
    memory[3173] = 32'h3e017d9b ;
    memory[3174] = 32'hbd27a8d4 ;
    memory[3175] = 32'hbda8aa24 ;
    memory[3176] = 32'h3cb1e788 ;
    memory[3177] = 32'h3e299eee ;
    memory[3178] = 32'hbdd907af ;
    memory[3179] = 32'hbd47d3b5 ;
    memory[3180] = 32'hbe0e5035 ;
    memory[3181] = 32'h3dc5d97d ;
    memory[3182] = 32'hbd1b0594 ;
    memory[3183] = 32'hbe420a6c ;
    memory[3184] = 32'hbdfdb561 ;
    memory[3185] = 32'h3d72329b ;
    memory[3186] = 32'h3d3e74d0 ;
    memory[3187] = 32'h3b9884c4 ;
    memory[3188] = 32'h3de2fdfe ;
    memory[3189] = 32'hbe21bf32 ;
    memory[3190] = 32'hbdd0a139 ;
    memory[3191] = 32'hbcf0ab03 ;
    memory[3192] = 32'h3dafd4ba ;
    memory[3193] = 32'hbdb624af ;
    memory[3194] = 32'h3e215520 ;
    memory[3195] = 32'h3dd4fe58 ;
    memory[3196] = 32'h3d1cdc6e ;
    memory[3197] = 32'h3e03b6d1 ;
    memory[3198] = 32'hbe1dc229 ;
    memory[3199] = 32'hbdd30395 ;
end



endmodule
